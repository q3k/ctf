module dut(input [39:0] lever, output lamp_1_1938);

assign lamp_1_1938 = gate3_1_1934;
assign gate3_1_1934 = gate3_1_1929 & gate3_4_1929;
assign gate3_4_1929 = gate3_7_1915 & not_5_1928;
assign not_5_1928 = ~gate3_4_1922;
assign gate3_4_1922 = gate3_1_1915 & not_5_1921;
assign not_5_1921 = ~gate3_4_1915;
assign gate3_4_1915 = gate3_1_1908 & gate3_100_1628;
assign gate3_100_1628 = xor_69_1576 & not_101_1627;
assign not_101_1627 = ~gate3_93_1602;
assign gate3_93_1602 = gate3_73_1576 & xor_82_1576;
assign xor_82_1576 = gate3_84_1555 ^ not_113_1529;
assign not_113_1529 = ~xor_113_1528;
assign xor_113_1528 = gate3_80_728 ^ not_85_1504;
assign not_85_1504 = ~xor_85_1503;
assign xor_85_1503 = not_114_1454 ^ gate3_92_1478;
assign gate3_92_1478 = gate3_88_1430 & gate3_100_1453;
assign gate3_100_1453 = gate3_179_1394 | xor_167_1430;
assign xor_167_1430 = gate3_168_1394 ^ not_182_1395;
assign not_182_1395 = ~xor_182_1394;
assign xor_182_1394 = not_187_1367 ^ xor_391_774;
assign xor_391_774 = gate3_440_728 ^ gate3_452_728;
assign gate3_452_728 = lever[34] & lever[18];
assign gate3_440_728 = lever[19] & lever[33];
assign not_187_1367 = ~xor_187_1366;
assign xor_187_1366 = gate3_188_1330 ^ xor_191_1330;
assign xor_191_1330 = gate3_229_1108 ^ not_201_1280;
assign not_201_1280 = ~xor_201_1279;
assign xor_201_1279 = not_216_1234 ^ gate3_446_728;
assign gate3_446_728 = lever[14] & lever[38];
assign not_216_1234 = ~xor_216_1233;
assign xor_216_1233 = xor_241_1108 ^ gate3_182_1182;
assign gate3_182_1182 = gate3_239_1054 | gate3_220_1108;
assign gate3_220_1108 = not_221_1107 & gate3_198_983;
assign gate3_198_983 = gate3_340_774 | gate3_291_857;
assign gate3_291_857 = gate3_404_728 & xor_343_774;
assign xor_343_774 = gate3_329_728 ^ gate3_407_728;
assign gate3_407_728 = lever[15] & lever[35];
assign gate3_329_728 = lever[36] & lever[14];
assign gate3_404_728 = lever[13] & lever[37];
assign gate3_340_774 = gate3_329_728 & gate3_407_728;
assign not_221_1107 = ~xor_248_1054;
assign xor_248_1054 = not_315_858 ^ gate3_201_983;
assign gate3_201_983 = gate3_352_774 | gate3_300_857;
assign gate3_300_857 = gate3_413_728 & xor_355_774;
assign xor_355_774 = gate3_392_728 ^ gate3_416_728;
assign gate3_416_728 = lever[32] & lever[18];
assign gate3_392_728 = lever[17] & lever[33];
assign gate3_413_728 = lever[34] & lever[16];
assign gate3_352_774 = gate3_389_728 & gate3_419_728;
assign gate3_419_728 = lever[18] & lever[33];
assign gate3_389_728 = lever[32] & lever[17];
assign not_315_858 = ~xor_315_857;
assign xor_315_857 = xor_373_774 ^ gate3_425_728;
assign gate3_425_728 = lever[14] & lever[37];
assign xor_373_774 = gate3_410_728 ^ gate3_428_728;
assign gate3_428_728 = lever[35] & lever[16];
assign gate3_410_728 = lever[36] & lever[15];
assign gate3_239_1054 = gate3_201_983 & not_240_1053;
assign not_240_1053 = ~not_315_858;
assign xor_241_1108 = gate3_207_983 ^ xor_256_1054;
assign xor_256_1054 = not_325_858 ^ gate3_210_983;
assign gate3_210_983 = gate3_376_774 | gate3_318_857;
assign gate3_318_857 = gate3_434_728 & xor_379_774;
assign xor_379_774 = gate3_419_728 ^ gate3_437_728;
assign gate3_437_728 = lever[32] & lever[19];
assign gate3_434_728 = lever[17] & lever[34];
assign gate3_376_774 = gate3_416_728 & gate3_440_728;
assign not_325_858 = ~xor_325_857;
assign xor_325_857 = gate3_449_728 ^ xor_388_774;
assign xor_388_774 = gate3_431_728 ^ gate3_95_728;
assign gate3_95_728 = lever[35] & lever[17];
assign gate3_431_728 = lever[16] & lever[36];
assign gate3_449_728 = lever[15] & lever[37];
assign gate3_207_983 = gate3_370_774 | gate3_309_857;
assign gate3_309_857 = gate3_425_728 & xor_373_774;
assign gate3_370_774 = gate3_407_728 & gate3_431_728;
assign gate3_229_1108 = gate3_253_1054 | not_322_858;
assign not_322_858 = ~xor_322_857;
assign xor_322_857 = gate3_434_728 ^ xor_379_774;
assign gate3_253_1054 = gate3_288_857 & gate3_191_983;
assign gate3_191_983 = gate3_361_774 | not_303_858;
assign not_303_858 = ~xor_303_857;
assign xor_303_857 = gate3_413_728 ^ xor_355_774;
assign gate3_361_774 = gate3_359_728 | not_362_773;
assign not_362_773 = ~gate3_398_728;
assign gate3_398_728 = lever[19] & lever[31];
assign gate3_359_728 = lever[30] & lever[18];
assign gate3_288_857 = not_359_774 | not_289_856;
assign not_289_856 = ~gate3_398_728;
assign not_359_774 = ~gate3_359_728;
assign gate3_188_1330 = gate3_191_1279 | gate3_210_1233;
assign gate3_210_1233 = not_211_1232 & gate3_172_1182;
assign gate3_172_1182 = gate3_233_1054 | gate3_211_1108;
assign gate3_211_1108 = gate3_182_983 & not_212_1107;
assign not_212_1107 = ~xor_236_1054;
assign xor_236_1054 = not_297_858 ^ gate3_188_983;
assign gate3_188_983 = gate3_328_774 | gate3_276_857;
assign gate3_276_857 = gate3_386_728 & xor_331_774;
assign xor_331_774 = gate3_335_728 ^ gate3_389_728;
assign gate3_335_728 = lever[16] & lever[33];
assign gate3_386_728 = lever[34] & lever[15];
assign gate3_328_774 = gate3_335_728 & gate3_389_728;
assign not_297_858 = ~xor_297_857;
assign xor_297_857 = gate3_404_728 ^ xor_343_774;
assign gate3_182_983 = gate3_280_774 | gate3_231_857;
assign gate3_231_857 = gate3_323_728 & xor_283_774;
assign xor_283_774 = gate3_308_728 ^ gate3_326_728;
assign gate3_326_728 = lever[35] & lever[14];
assign gate3_308_728 = lever[13] & lever[36];
assign gate3_323_728 = lever[12] & lever[37];
assign gate3_280_774 = gate3_308_728 & gate3_326_728;
assign gate3_233_1054 = gate3_188_983 & not_234_1053;
assign not_234_1053 = ~not_297_858;
assign not_211_1232 = ~xor_223_1108;
assign xor_223_1108 = gate3_198_983 ^ xor_248_1054;
assign gate3_191_1279 = gate3_422_728 & not_213_1234;
assign not_213_1234 = ~xor_213_1233;
assign xor_213_1233 = gate3_172_1182 ^ xor_223_1108;
assign gate3_422_728 = lever[13] & lever[38];
assign gate3_168_1394 = not_184_1367 | not_169_1393;
assign not_169_1393 = ~xor_235_1108;
assign xor_235_1108 = gate3_253_1054 ^ not_322_858;
assign not_184_1367 = ~xor_184_1366;
assign xor_184_1366 = gate3_179_1330 ^ not_185_1331;
assign not_185_1331 = ~xor_185_1330;
assign xor_185_1330 = gate3_204_1233 ^ not_198_1280;
assign not_198_1280 = ~xor_198_1279;
assign xor_198_1279 = gate3_422_728 ^ not_213_1234;
assign gate3_204_1233 = gate3_164_1182 | not_205_1232;
assign not_205_1232 = ~xor_194_983;
assign xor_194_983 = not_303_858 ^ gate3_361_774;
assign gate3_164_1182 = gate3_227_1054 & gate3_196_1108;
assign gate3_196_1108 = not_282_858 | xor_230_1054;
assign xor_230_1054 = gate3_176_983 ^ not_334_775;
assign not_334_775 = ~xor_334_774;
assign xor_334_774 = gate3_374_728 ^ gate3_395_728;
assign gate3_395_728 = lever[31] & lever[18];
assign gate3_374_728 = lever[30] & lever[19];
assign gate3_176_983 = gate3_307_774 | gate3_256_857;
assign gate3_256_857 = gate3_368_728 & xor_310_774;
assign xor_310_774 = gate3_371_728 ^ gate3_359_728;
assign gate3_371_728 = lever[29] & lever[19];
assign gate3_368_728 = lever[31] & lever[17];
assign gate3_307_774 = gate3_356_728 & gate3_374_728;
assign gate3_356_728 = lever[29] & lever[18];
assign not_282_858 = ~xor_282_857;
assign xor_282_857 = gate3_386_728 ^ xor_331_774;
assign gate3_227_1054 = not_334_775 | not_228_1053;
assign not_228_1053 = ~gate3_176_983;
assign gate3_179_1330 = gate3_196_1233 & not_180_1329;
assign not_180_1329 = ~gate3_185_1279;
assign gate3_185_1279 = gate3_401_728 & not_201_1234;
assign not_201_1234 = ~xor_201_1233;
assign xor_201_1233 = xor_214_1108 ^ gate3_151_1182;
assign gate3_151_1182 = gate3_164_1108 | gate3_200_1054;
assign gate3_200_1054 = gate3_162_983 & not_201_1053;
assign not_201_1053 = ~not_237_858;
assign not_237_858 = ~xor_237_857;
assign xor_237_857 = gate3_323_728 ^ xor_283_774;
assign gate3_162_983 = gate3_286_774 | gate3_240_857;
assign gate3_240_857 = gate3_338_728 & xor_292_774;
assign xor_292_774 = gate3_314_728 ^ gate3_332_728;
assign gate3_332_728 = lever[32] & lever[16];
assign gate3_314_728 = lever[15] & lever[33];
assign gate3_338_728 = lever[14] & lever[34];
assign gate3_286_774 = gate3_314_728 & gate3_332_728;
assign gate3_164_1108 = gate3_158_983 & not_165_1107;
assign not_165_1107 = ~xor_205_1054;
assign xor_205_1054 = not_237_858 ^ gate3_162_983;
assign gate3_158_983 = gate3_268_774 | gate3_217_857;
assign gate3_217_857 = gate3_302_728 & xor_271_774;
assign xor_271_774 = gate3_275_728 ^ gate3_305_728;
assign gate3_305_728 = lever[13] & lever[35];
assign gate3_275_728 = lever[12] & lever[36];
assign gate3_302_728 = lever[11] & lever[37];
assign gate3_268_774 = gate3_275_728 & gate3_305_728;
assign xor_214_1108 = xor_236_1054 ^ gate3_182_983;
assign gate3_401_728 = lever[12] & lever[38];
assign gate3_196_1233 = not_197_1232 | xor_214_1108;
assign not_197_1232 = ~gate3_151_1182;
assign gate3_179_1394 = gate3_179_1366 & gate3_182_1330;
assign gate3_182_1330 = gate3_204_1233 | not_198_1280;
assign gate3_179_1366 = gate3_179_1330 | not_185_1331;
assign gate3_88_1430 = gate3_168_1394 | not_89_1429;
assign not_89_1429 = ~not_182_1395;
assign not_114_1454 = ~xor_114_1453;
assign xor_114_1453 = gate3_106_1394 ^ xor_111_1430;
assign xor_111_1430 = gate3_121_1394 ^ xor_114_1394;
assign xor_114_1394 = gate3_101_728 ^ xor_121_1366;
assign xor_121_1366 = not_111_1280 ^ gate3_95_1330;
assign gate3_95_1330 = gate3_117_1233 | gate3_97_1279;
assign gate3_97_1279 = gate3_446_728 & not_216_1234;
assign gate3_117_1233 = gate3_182_1182 & not_118_1232;
assign not_118_1232 = ~xor_241_1108;
assign not_111_1280 = ~xor_111_1279;
assign xor_111_1279 = gate3_83_728 ^ not_124_1234;
assign not_124_1234 = ~xor_124_1233;
assign xor_124_1233 = xor_115_1054 ^ gate3_51_1182;
assign gate3_51_1182 = gate3_109_1054 | gate3_95_1108;
assign gate3_95_1108 = gate3_207_983 & not_96_1107;
assign not_96_1107 = ~xor_256_1054;
assign gate3_109_1054 = gate3_210_983 & not_110_1053;
assign not_110_1053 = ~not_325_858;
assign xor_115_1054 = gate3_38_983 ^ xor_49_983;
assign xor_49_983 = gate3_112_774 ^ not_99_858;
assign not_99_858 = ~xor_99_857;
assign xor_99_857 = gate3_86_728 ^ xor_97_774;
assign xor_97_774 = gate3_98_728 ^ gate3_89_728;
assign gate3_89_728 = lever[18] & lever[35];
assign gate3_98_728 = lever[17] & lever[36];
assign gate3_86_728 = lever[37] & lever[16];
assign gate3_112_774 = gate3_419_728 & gate3_101_728;
assign gate3_101_728 = lever[34] & lever[19];
assign gate3_38_983 = gate3_91_774 | gate3_88_857;
assign gate3_88_857 = gate3_449_728 & xor_388_774;
assign gate3_91_774 = gate3_431_728 & gate3_95_728;
assign gate3_83_728 = lever[15] & lever[38];
assign gate3_121_1394 = not_187_1367 | not_122_1393;
assign not_122_1393 = ~xor_391_774;
assign gate3_106_1394 = gate3_91_1330 & not_107_1393;
assign not_107_1393 = ~gate3_111_1366;
assign gate3_111_1366 = xor_191_1330 & gate3_188_1330;
assign gate3_91_1330 = gate3_229_1108 | not_201_1280;
assign gate3_80_728 = lever[14] & lever[39];
assign gate3_84_1555 = gate3_67_1503 | gate3_100_1528;
assign gate3_100_1528 = gate3_443_728 & not_121_1504;
assign not_121_1504 = ~xor_121_1503;
assign xor_121_1503 = gate3_137_1478 ^ xor_170_1453;
assign xor_170_1453 = gate3_179_1394 ^ xor_167_1430;
assign gate3_137_1478 = gate3_159_1430 & gate3_164_1453;
assign gate3_164_1453 = gate3_165_1394 | not_162_1431;
assign not_162_1431 = ~xor_162_1430;
assign xor_162_1430 = xor_171_1394 ^ gate3_159_1394;
assign gate3_159_1394 = not_160_1393 | xor_172_1366;
assign xor_172_1366 = xor_170_1330 ^ gate3_159_1330;
assign gate3_159_1330 = not_160_1329 & gate3_170_1233;
assign gate3_170_1233 = xor_170_1108 | not_171_1232;
assign not_171_1232 = ~gate3_139_1182;
assign gate3_139_1182 = gate3_190_1054 | gate3_151_1108;
assign gate3_151_1108 = not_152_1107 & gate3_139_983;
assign gate3_139_983 = gate3_229_774 | gate3_199_857;
assign gate3_199_857 = gate3_263_728 & xor_232_774;
assign xor_232_774 = gate3_269_728 ^ gate3_266_728;
assign gate3_266_728 = lever[36] & lever[11];
assign gate3_269_728 = lever[12] & lever[35];
assign gate3_263_728 = lever[10] & lever[37];
assign gate3_229_774 = gate3_266_728 & gate3_269_728;
assign not_152_1107 = ~xor_196_1054;
assign xor_196_1054 = not_223_858 ^ gate3_145_983;
assign gate3_145_983 = gate3_274_774 | gate3_226_857;
assign gate3_226_857 = gate3_317_728 & xor_277_774;
assign xor_277_774 = gate3_311_728 ^ gate3_284_728;
assign gate3_284_728 = lever[14] & lever[33];
assign gate3_311_728 = lever[32] & lever[15];
assign gate3_317_728 = lever[34] & lever[13];
assign gate3_274_774 = gate3_284_728 & gate3_311_728;
assign not_223_858 = ~xor_223_857;
assign xor_223_857 = gate3_302_728 ^ xor_271_774;
assign gate3_190_1054 = gate3_145_983 & not_191_1053;
assign not_191_1053 = ~not_223_858;
assign xor_170_1108 = xor_205_1054 ^ gate3_158_983;
assign not_160_1329 = ~gate3_172_1279;
assign gate3_172_1279 = gate3_320_728 & not_182_1234;
assign not_182_1234 = ~xor_182_1233;
assign xor_182_1233 = gate3_139_1182 ^ xor_170_1108;
assign gate3_320_728 = lever[11] & lever[38];
assign xor_170_1330 = gate3_193_1233 ^ not_188_1280;
assign not_188_1280 = ~xor_188_1279;
assign xor_188_1279 = gate3_401_728 ^ not_201_1234;
assign gate3_193_1233 = gate3_148_1182 | not_194_1232;
assign not_194_1232 = ~xor_205_1108;
assign xor_205_1108 = not_282_858 ^ xor_230_1054;
assign gate3_148_1182 = gate3_209_1054 & gate3_182_1108;
assign gate3_182_1108 = xor_212_1054 | not_246_858;
assign not_246_858 = ~xor_246_857;
assign xor_246_857 = gate3_338_728 ^ xor_292_774;
assign xor_212_1054 = not_259_858 ^ gate3_165_983;
assign gate3_165_983 = gate3_295_774 | gate3_252_857;
assign gate3_252_857 = gate3_365_728 & xor_304_774;
assign xor_304_774 = gate3_353_728 ^ gate3_356_728;
assign gate3_353_728 = lever[30] & lever[17];
assign gate3_365_728 = lever[16] & lever[31];
assign gate3_295_774 = gate3_359_728 & gate3_362_728;
assign gate3_362_728 = lever[29] & lever[17];
assign not_259_858 = ~xor_259_857;
assign xor_259_857 = gate3_368_728 ^ xor_310_774;
assign gate3_209_1054 = not_259_858 | not_210_1053;
assign not_210_1053 = ~gate3_165_983;
assign not_160_1393 = ~not_207_1234;
assign not_207_1234 = ~xor_207_1233;
assign xor_207_1233 = gate3_164_1182 ^ xor_194_983;
assign xor_171_1394 = not_184_1367 ^ xor_235_1108;
assign gate3_165_1394 = gate3_164_1330 & gate3_169_1366;
assign gate3_169_1366 = gate3_159_1330 | not_170_1365;
assign not_170_1365 = ~xor_170_1330;
assign gate3_164_1330 = gate3_193_1233 | not_188_1280;
assign gate3_159_1430 = gate3_159_1394 | xor_171_1394;
assign gate3_443_728 = lever[13] & lever[39];
assign gate3_67_1503 = xor_170_1453 & not_68_1502;
assign not_68_1502 = ~gate3_137_1478;
assign gate3_73_1576 = not_97_1529 | not_74_1575;
assign not_74_1575 = ~gate3_81_1555;
assign gate3_81_1555 = gate3_116_1503 | gate3_151_1528;
assign gate3_151_1528 = gate3_77_728 & not_57_1504;
assign not_57_1504 = ~xor_57_1503;
assign xor_57_1503 = gate3_134_1478 ^ xor_167_1453;
assign xor_167_1453 = not_162_1431 ^ gate3_165_1394;
assign gate3_134_1478 = gate3_161_1453 & gate3_156_1430;
assign gate3_156_1430 = xor_162_1394 | gate3_156_1394;
assign gate3_156_1394 = not_106_1367 | not_157_1393;
assign not_157_1393 = ~not_114_1234;
assign not_114_1234 = ~xor_114_1233;
assign xor_114_1233 = gate3_148_1182 ^ xor_205_1108;
assign not_106_1367 = ~xor_106_1366;
assign xor_106_1366 = gate3_139_1330 ^ not_156_1331;
assign not_156_1331 = ~xor_156_1330;
assign xor_156_1330 = gate3_182_1279 ^ not_179_1280;
assign not_179_1280 = ~xor_179_1279;
assign xor_179_1279 = gate3_320_728 ^ not_182_1234;
assign gate3_182_1279 = gate3_185_1233 & gate3_145_1182;
assign gate3_145_1182 = gate3_243_857 | not_146_1181;
assign not_146_1181 = ~xor_186_1108;
assign xor_186_1108 = not_246_858 ^ xor_212_1054;
assign gate3_243_857 = not_347_774 | not_244_856;
assign not_244_856 = ~gate3_350_728;
assign gate3_350_728 = lever[28] & lever[19];
assign not_347_774 = ~gate3_347_728;
assign gate3_347_728 = lever[27] & lever[18];
assign gate3_185_1233 = gate3_35_1182 | xor_47_1182;
assign xor_47_1182 = gate3_243_857 ^ xor_186_1108;
assign gate3_35_1182 = gate3_218_1054 & gate3_192_1108;
assign gate3_192_1108 = not_270_858 | xor_221_1054;
assign xor_221_1054 = gate3_168_983 ^ not_265_858;
assign not_265_858 = ~xor_265_857;
assign xor_265_857 = gate3_365_728 ^ xor_304_774;
assign gate3_168_983 = gate3_313_774 | gate3_262_857;
assign gate3_262_857 = gate3_383_728 & xor_325_774;
assign xor_325_774 = gate3_362_728 ^ gate3_377_728;
assign gate3_377_728 = lever[30] & lever[16];
assign gate3_383_728 = lever[31] & lever[15];
assign gate3_313_774 = gate3_362_728 & gate3_377_728;
assign not_270_858 = ~xor_270_857;
assign xor_270_857 = gate3_317_728 ^ xor_277_774;
assign gate3_218_1054 = not_265_858 | not_219_1053;
assign not_219_1053 = ~gate3_168_983;
assign gate3_139_1330 = gate3_164_1233 & not_140_1329;
assign not_140_1329 = ~gate3_166_1279;
assign gate3_166_1279 = gate3_68_728 & xor_97_1233;
assign xor_97_1233 = gate3_133_1182 ^ xor_158_1108;
assign xor_158_1108 = gate3_139_983 ^ xor_196_1054;
assign gate3_133_1182 = gate3_148_1108 & gate3_184_1054;
assign gate3_184_1054 = not_205_858 | not_185_1053;
assign not_185_1053 = ~gate3_124_983;
assign gate3_124_983 = gate3_208_857 | gate3_235_774;
assign gate3_235_774 = gate3_278_728 & gate3_281_728;
assign gate3_281_728 = lever[13] & lever[33];
assign gate3_278_728 = lever[32] & lever[14];
assign gate3_208_857 = gate3_290_728 & xor_238_774;
assign xor_238_774 = gate3_278_728 ^ gate3_281_728;
assign gate3_290_728 = lever[12] & lever[34];
assign not_205_858 = ~xor_205_857;
assign xor_205_857 = gate3_263_728 ^ xor_232_774;
assign gate3_148_1108 = xor_187_1054 | not_149_1107;
assign not_149_1107 = ~gate3_129_983;
assign gate3_129_983 = gate3_250_774 | gate3_213_857;
assign gate3_213_857 = gate3_299_728 & xor_265_774;
assign xor_265_774 = gate3_272_728 ^ gate3_293_728;
assign gate3_293_728 = lever[36] & lever[10];
assign gate3_272_728 = lever[11] & lever[35];
assign gate3_299_728 = lever[9] & lever[37];
assign gate3_250_774 = gate3_272_728 & gate3_293_728;
assign xor_187_1054 = not_205_858 ^ gate3_124_983;
assign gate3_68_728 = lever[10] & lever[38];
assign gate3_164_1233 = gate3_133_1182 | xor_158_1108;
assign xor_162_1394 = xor_172_1366 ^ not_207_1234;
assign gate3_161_1453 = gate3_101_1394 | not_85_1431;
assign not_85_1431 = ~xor_85_1430;
assign xor_85_1430 = gate3_156_1394 ^ xor_162_1394;
assign gate3_101_1394 = gate3_145_1330 & gate3_166_1366;
assign gate3_166_1366 = gate3_139_1330 | not_156_1331;
assign gate3_145_1330 = not_179_1280 | gate3_182_1279;
assign gate3_77_728 = lever[12] & lever[39];
assign gate3_116_1503 = xor_167_1453 & not_117_1502;
assign not_117_1502 = ~gate3_134_1478;
assign not_97_1529 = ~xor_97_1528;
assign xor_97_1528 = gate3_443_728 ^ not_121_1504;
assign xor_69_1576 = gate3_81_1555 ^ not_97_1529;
assign gate3_1_1908 = gate3_1_1901 & gate3_67_1654;
assign gate3_67_1654 = gate3_75_1602 & gate3_95_1628;
assign gate3_95_1628 = xor_84_1602 | gate3_87_1602;
assign gate3_87_1602 = not_77_1556 | not_88_1601;
assign not_88_1601 = ~gate3_66_1576;
assign gate3_66_1576 = gate3_79_1528 | gate3_67_1555;
assign gate3_67_1555 = gate3_71_728 & not_84_1529;
assign not_84_1529 = ~xor_84_1528;
assign xor_84_1528 = xor_87_1478 ^ gate3_51_1503;
assign gate3_51_1503 = gate3_54_1478 & gate3_82_1453;
assign gate3_82_1453 = not_90_1395 | gate3_67_1430;
assign gate3_67_1430 = gate3_67_1394 & gate3_82_1366;
assign gate3_82_1366 = gate3_232_1330 | not_301_1280;
assign not_301_1280 = ~xor_301_1279;
assign xor_301_1279 = xor_294_1233 ^ gate3_619_774;
assign gate3_619_774 = gate3_350_728 & not_620_773;
assign not_620_773 = ~gate3_347_728;
assign xor_294_1233 = gate3_265_1182 ^ xor_268_1182;
assign xor_268_1182 = xor_354_1108 ^ gate3_346_1108;
assign gate3_346_1108 = not_347_1107 | not_317_1054;
assign not_317_1054 = ~gate3_317_983;
assign gate3_317_983 = gate3_607_774 | gate3_513_857;
assign gate3_513_857 = gate3_680_728 & xor_613_774;
assign xor_613_774 = gate3_683_728 ^ gate3_347_728;
assign gate3_683_728 = lever[26] & lever[19];
assign gate3_680_728 = lever[28] & lever[17];
assign gate3_607_774 = gate3_341_728 & gate3_608_728;
assign gate3_608_728 = lever[26] & lever[18];
assign gate3_341_728 = lever[27] & lever[19];
assign not_347_1107 = ~xor_616_774;
assign xor_616_774 = gate3_344_728 ^ gate3_341_728;
assign gate3_344_728 = lever[28] & lever[18];
assign xor_354_1108 = not_270_858 ^ xor_221_1054;
assign gate3_265_1182 = gate3_339_1108 & gate3_376_1054;
assign gate3_376_1054 = not_531_858 | not_377_1053;
assign not_377_1053 = ~gate3_311_983;
assign gate3_311_983 = gate3_598_774 | gate3_504_857;
assign gate3_504_857 = gate3_677_728 & xor_601_774;
assign xor_601_774 = gate3_602_728 ^ gate3_380_728;
assign gate3_380_728 = lever[16] & lever[29];
assign gate3_602_728 = lever[15] & lever[30];
assign gate3_677_728 = lever[31] & lever[14];
assign gate3_598_774 = gate3_380_728 & gate3_602_728;
assign not_531_858 = ~xor_531_857;
assign xor_531_857 = gate3_383_728 ^ xor_325_774;
assign gate3_339_1108 = not_525_858 | xor_379_1054;
assign xor_379_1054 = gate3_311_983 ^ not_531_858;
assign not_525_858 = ~xor_525_857;
assign xor_525_857 = gate3_290_728 ^ xor_238_774;
assign gate3_232_1330 = not_288_1279 | not_382_1055;
assign not_382_1055 = ~xor_382_1054;
assign xor_382_1054 = gate3_317_983 ^ xor_616_774;
assign not_288_1279 = ~not_288_1234;
assign not_288_1234 = ~xor_288_1233;
assign xor_288_1233 = gate3_250_1182 ^ not_256_1183;
assign not_256_1183 = ~xor_256_1182;
assign xor_256_1182 = gate3_361_1054 ^ xor_343_1108;
assign xor_343_1108 = not_525_858 ^ xor_379_1054;
assign gate3_361_1054 = not_362_1053 | not_516_858;
assign not_516_858 = ~xor_516_857;
assign xor_516_857 = gate3_680_728 ^ xor_613_774;
assign not_362_1053 = ~gate3_302_983;
assign gate3_302_983 = gate3_529_774 | gate3_432_857;
assign gate3_432_857 = gate3_605_728 & xor_532_774;
assign xor_532_774 = gate3_521_728 ^ gate3_608_728;
assign gate3_521_728 = lever[27] & lever[17];
assign gate3_605_728 = lever[28] & lever[16];
assign gate3_529_774 = gate3_347_728 & gate3_518_728;
assign gate3_518_728 = lever[26] & lever[17];
assign gate3_250_1182 = gate3_352_1054 & gate3_318_1108;
assign gate3_318_1108 = not_501_858 | xor_355_1054;
assign xor_355_1054 = gate3_299_983 ^ not_507_858;
assign not_507_858 = ~xor_507_857;
assign xor_507_857 = gate3_677_728 ^ xor_601_774;
assign gate3_299_983 = gate3_520_774 | gate3_424_857;
assign gate3_424_857 = gate3_596_728 & xor_523_774;
assign xor_523_774 = gate3_599_728 ^ gate3_584_728;
assign gate3_584_728 = lever[14] & lever[30];
assign gate3_599_728 = lever[29] & lever[15];
assign gate3_596_728 = lever[31] & lever[13];
assign gate3_520_774 = gate3_584_728 & gate3_599_728;
assign not_501_858 = ~xor_501_857;
assign xor_501_857 = gate3_674_728 ^ xor_592_774;
assign xor_592_774 = gate3_287_728 ^ gate3_593_728;
assign gate3_593_728 = lever[12] & lever[33];
assign gate3_287_728 = lever[32] & lever[13];
assign gate3_674_728 = lever[11] & lever[34];
assign gate3_352_1054 = not_507_858 | not_353_1053;
assign not_353_1053 = ~gate3_299_983;
assign gate3_67_1394 = not_231_1367 | not_68_1393;
assign not_68_1393 = ~xor_237_1366;
assign xor_237_1366 = not_301_1280 ^ gate3_232_1330;
assign not_231_1367 = ~xor_231_1366;
assign xor_231_1366 = gate3_237_1330 ^ not_243_1331;
assign not_243_1331 = ~xor_243_1330;
assign xor_243_1330 = gate3_296_1279 ^ not_293_1280;
assign not_293_1280 = ~xor_293_1279;
assign xor_293_1279 = gate3_695_728 ^ xor_291_1233;
assign xor_291_1233 = gate3_262_1182 ^ xor_349_1108;
assign xor_349_1108 = gate3_129_983 ^ xor_187_1054;
assign gate3_262_1182 = gate3_370_1054 & gate3_329_1108;
assign gate3_329_1108 = xor_373_1054 | not_330_1107;
assign not_330_1107 = ~gate3_305_983;
assign gate3_305_983 = gate3_580_774 | gate3_483_857;
assign gate3_483_857 = gate3_671_728 & xor_583_774;
assign xor_583_774 = gate3_296_728 ^ gate3_665_728;
assign gate3_665_728 = lever[36] & lever[9];
assign gate3_296_728 = lever[35] & lever[10];
assign gate3_671_728 = lever[8] & lever[37];
assign gate3_580_774 = gate3_665_728 & gate3_296_728;
assign xor_373_1054 = not_522_858 ^ gate3_308_983;
assign gate3_308_983 = gate3_589_774 | gate3_495_857;
assign gate3_495_857 = gate3_674_728 & xor_592_774;
assign gate3_589_774 = gate3_590_728 & gate3_281_728;
assign gate3_590_728 = lever[32] & lever[12];
assign not_522_858 = ~xor_522_857;
assign xor_522_857 = gate3_299_728 ^ xor_265_774;
assign gate3_370_1054 = not_522_858 | not_371_1053;
assign not_371_1053 = ~gate3_308_983;
assign gate3_695_728 = lever[9] & lever[38];
assign gate3_296_1279 = gate3_253_1182 & gate3_283_1233;
assign gate3_283_1233 = gate3_250_1182 | not_284_1232;
assign not_284_1232 = ~not_256_1183;
assign gate3_253_1182 = gate3_361_1054 | not_254_1181;
assign not_254_1181 = ~xor_343_1108;
assign gate3_237_1330 = not_238_1329 & gate3_273_1233;
assign gate3_273_1233 = gate3_247_1182 | xor_336_1108;
assign xor_336_1108 = gate3_305_983 ^ xor_373_1054;
assign gate3_247_1182 = gate3_341_1054 & gate3_309_1108;
assign gate3_309_1108 = xor_344_1054 | not_310_1107;
assign not_310_1107 = ~gate3_290_983;
assign gate3_290_983 = gate3_571_774 | gate3_474_857;
assign gate3_474_857 = gate3_659_728 & xor_574_774;
assign xor_574_774 = gate3_650_728 ^ gate3_662_728;
assign gate3_662_728 = lever[9] & lever[35];
assign gate3_650_728 = lever[36] & lever[8];
assign gate3_659_728 = lever[7] & lever[37];
assign gate3_571_774 = gate3_650_728 & gate3_662_728;
assign xor_344_1054 = not_489_858 ^ gate3_293_983;
assign gate3_293_983 = gate3_511_774 | gate3_417_857;
assign gate3_417_857 = gate3_587_728 & xor_517_774;
assign xor_517_774 = gate3_575_728 ^ gate3_590_728;
assign gate3_575_728 = lever[33] & lever[11];
assign gate3_587_728 = lever[10] & lever[34];
assign gate3_511_774 = gate3_575_728 & gate3_590_728;
assign not_489_858 = ~xor_489_857;
assign xor_489_857 = gate3_671_728 ^ xor_583_774;
assign gate3_341_1054 = not_489_858 | not_342_1053;
assign not_342_1053 = ~gate3_293_983;
assign not_238_1329 = ~gate3_280_1279;
assign gate3_280_1279 = gate3_686_728 & xor_277_1233;
assign xor_277_1233 = gate3_247_1182 ^ xor_336_1108;
assign gate3_686_728 = lever[8] & lever[38];
assign not_90_1395 = ~xor_90_1394;
assign xor_90_1394 = not_88_1331 ^ not_98_1367;
assign not_98_1367 = ~xor_98_1366;
assign xor_98_1366 = gate3_57_1330 ^ not_82_1331;
assign not_82_1331 = ~xor_82_1330;
assign xor_82_1330 = not_67_1280 ^ gate3_82_1279;
assign gate3_82_1279 = gate3_26_1182 & gate3_106_1233;
assign gate3_106_1233 = xor_268_1182 | gate3_265_1182;
assign gate3_26_1182 = gate3_346_1108 | not_27_1181;
assign not_27_1181 = ~xor_354_1108;
assign not_67_1280 = ~xor_67_1279;
assign xor_67_1279 = gate3_68_728 ^ xor_97_1233;
assign gate3_57_1330 = not_58_1329 & gate3_88_1233;
assign gate3_88_1233 = gate3_262_1182 | xor_349_1108;
assign not_58_1329 = ~gate3_56_1279;
assign gate3_56_1279 = gate3_695_728 & xor_291_1233;
assign not_88_1331 = ~xor_88_1330;
assign xor_88_1330 = gate3_90_1279 ^ xor_109_1233;
assign xor_109_1233 = gate3_35_1182 ^ xor_47_1182;
assign gate3_90_1279 = xor_294_1233 & gate3_619_774;
assign gate3_54_1478 = gate3_53_1394 | not_55_1477;
assign not_55_1477 = ~xor_85_1453;
assign xor_85_1453 = gate3_67_1430 ^ not_90_1395;
assign gate3_53_1394 = gate3_54_1330 & gate3_69_1366;
assign gate3_69_1366 = gate3_237_1330 | not_243_1331;
assign gate3_54_1330 = not_293_1280 | gate3_296_1279;
assign xor_87_1478 = gate3_95_1394 ^ xor_93_1453;
assign xor_93_1453 = gate3_82_1430 ^ xor_98_1394;
assign xor_98_1394 = not_106_1367 ^ not_114_1234;
assign gate3_82_1430 = not_83_1429 | gate3_85_1330;
assign gate3_85_1330 = gate3_90_1279 & xor_109_1233;
assign not_83_1429 = ~gate3_87_1394;
assign gate3_87_1394 = not_88_1331 | not_98_1367;
assign gate3_95_1394 = gate3_67_1330 & gate3_95_1366;
assign gate3_95_1366 = gate3_57_1330 | not_82_1331;
assign gate3_67_1330 = not_67_1280 | gate3_82_1279;
assign gate3_71_728 = lever[10] & lever[39];
assign gate3_79_1528 = xor_87_1478 & not_80_1527;
assign not_80_1527 = ~gate3_51_1503;
assign not_77_1556 = ~xor_77_1555;
assign xor_77_1555 = not_91_1529 ^ gate3_74_728;
assign gate3_74_728 = lever[39] & lever[11];
assign not_91_1529 = ~xor_91_1528;
assign xor_91_1528 = xor_97_1453 ^ gate3_54_1503;
assign gate3_54_1503 = gate3_84_1478 & gate3_90_1453;
assign gate3_90_1453 = xor_98_1394 | not_91_1452;
assign not_91_1452 = ~gate3_82_1430;
assign gate3_84_1478 = gate3_95_1394 | xor_93_1453;
assign xor_97_1453 = gate3_101_1394 ^ not_85_1431;
assign xor_84_1602 = not_94_1529 ^ gate3_57_1576;
assign gate3_57_1576 = gate3_87_1528 | gate3_74_1555;
assign gate3_74_1555 = gate3_74_728 & not_91_1529;
assign gate3_87_1528 = xor_97_1453 & not_88_1527;
assign not_88_1527 = ~gate3_54_1503;
assign not_94_1529 = ~xor_94_1528;
assign xor_94_1528 = gate3_77_728 ^ not_57_1504;
assign gate3_75_1602 = not_94_1529 | not_76_1601;
assign not_76_1601 = ~gate3_57_1576;
assign gate3_1_1901 = gate3_92_1628 | gate3_1_1892;
assign gate3_1_1892 = gate3_1_1885 & gate3_127_1679;
assign gate3_127_1679 = gate3_71_1602 & gate3_64_1654;
assign gate3_64_1654 = gate3_66_1602 | gate3_77_1628;
assign gate3_77_1628 = not_64_1556 | not_78_1627;
assign not_78_1627 = ~gate3_57_1602;
assign gate3_57_1602 = gate3_49_1555 | gate3_51_1576;
assign gate3_51_1576 = gate3_692_728 & not_142_1556;
assign not_142_1556 = ~xor_142_1555;
assign xor_142_1555 = not_162_1479 ^ gate3_157_1528;
assign gate3_157_1528 = gate3_156_1478 & gate3_131_1503;
assign gate3_131_1503 = gate3_190_1430 | not_132_1502;
assign not_132_1502 = ~xor_159_1478;
assign xor_159_1478 = gate3_179_1453 ^ not_216_1395;
assign not_216_1395 = ~xor_216_1394;
assign xor_216_1394 = not_219_1367 ^ xor_228_1366;
assign xor_228_1366 = gate3_229_1330 ^ xor_290_1279;
assign xor_290_1279 = not_288_1234 ^ not_382_1055;
assign gate3_229_1330 = gate3_237_1182 | gate3_269_1279;
assign gate3_269_1279 = not_270_1234 & not_243_1183;
assign not_243_1183 = ~xor_243_1182;
assign xor_243_1182 = gate3_282_1108 ^ xor_364_1054;
assign xor_364_1054 = gate3_302_983 ^ not_516_858;
assign gate3_282_1108 = gate3_527_728 & not_283_1107;
assign not_283_1107 = ~xor_310_1054;
assign xor_310_1054 = gate3_248_983 ^ xor_256_983;
assign xor_256_983 = gate3_457_774 ^ not_438_858;
assign not_438_858 = ~xor_438_857;
assign xor_438_857 = gate3_605_728 ^ xor_532_774;
assign gate3_457_774 = gate3_476_728 & gate3_527_728;
assign gate3_527_728 = lever[25] & lever[19];
assign gate3_476_728 = lever[24] & lever[18];
assign gate3_248_983 = gate3_451_774 | gate3_366_857;
assign gate3_366_857 = xor_454_774 & gate3_515_728;
assign gate3_515_728 = lever[28] & lever[15];
assign xor_454_774 = gate3_512_728 ^ gate3_518_728;
assign gate3_512_728 = lever[27] & lever[16];
assign gate3_451_774 = gate3_512_728 & gate3_518_728;
assign not_270_1234 = ~xor_270_1233;
assign xor_270_1233 = gate3_219_1182 ^ xor_231_1182;
assign xor_231_1182 = xor_322_1108 ^ gate3_325_1108;
assign gate3_325_1108 = gate3_251_983 | gate3_307_1054;
assign gate3_307_1054 = gate3_248_983 & not_308_1053;
assign not_308_1053 = ~xor_256_983;
assign gate3_251_983 = gate3_457_774 & not_252_982;
assign not_252_982 = ~not_438_858;
assign xor_322_1108 = xor_355_1054 ^ not_501_858;
assign gate3_219_1182 = gate3_298_1054 & gate3_276_1108;
assign gate3_276_1108 = not_420_858 | xor_301_1054;
assign xor_301_1054 = not_429_858 ^ gate3_239_983;
assign gate3_239_983 = gate3_499_774 | gate3_408_857;
assign gate3_408_857 = gate3_578_728 & xor_508_774;
assign xor_508_774 = gate3_551_728 ^ gate3_581_728;
assign gate3_581_728 = lever[29] & lever[14];
assign gate3_551_728 = lever[13] & lever[30];
assign gate3_578_728 = lever[31] & lever[12];
assign gate3_499_774 = gate3_551_728 & gate3_581_728;
assign not_429_858 = ~xor_429_857;
assign xor_429_857 = gate3_596_728 ^ xor_523_774;
assign not_420_858 = ~xor_420_857;
assign xor_420_857 = gate3_587_728 ^ xor_517_774;
assign gate3_298_1054 = not_429_858 | not_299_1053;
assign not_299_1053 = ~gate3_239_983;
assign gate3_237_1182 = not_238_1181 & gate3_282_1108;
assign not_238_1181 = ~xor_364_1054;
assign not_219_1367 = ~xor_219_1366;
assign xor_219_1366 = gate3_220_1330 ^ xor_226_1330;
assign xor_226_1330 = not_283_1280 ^ gate3_286_1279;
assign gate3_286_1279 = gate3_225_1182 | gate3_267_1233;
assign gate3_267_1233 = xor_231_1182 & not_268_1232;
assign not_268_1232 = ~gate3_219_1182;
assign gate3_225_1182 = gate3_325_1108 & xor_322_1108;
assign not_283_1280 = ~xor_283_1279;
assign xor_283_1279 = gate3_686_728 ^ xor_277_1233;
assign gate3_220_1330 = gate3_261_1233 & not_221_1329;
assign not_221_1329 = ~gate3_263_1279;
assign gate3_263_1279 = not_264_1234 & gate3_668_728;
assign gate3_668_728 = lever[7] & lever[38];
assign not_264_1234 = ~xor_264_1233;
assign xor_264_1233 = gate3_216_1182 ^ xor_315_1108;
assign xor_315_1108 = gate3_290_983 ^ xor_344_1054;
assign gate3_216_1182 = gate3_334_1054 | gate3_303_1108;
assign gate3_303_1108 = not_304_1107 & gate3_278_983;
assign gate3_278_983 = gate3_562_774 | gate3_462_857;
assign gate3_462_857 = xor_565_774 & gate3_644_728;
assign gate3_644_728 = lever[6] & lever[37];
assign xor_565_774 = gate3_620_728 ^ gate3_647_728;
assign gate3_647_728 = lever[8] & lever[35];
assign gate3_620_728 = lever[7] & lever[36];
assign gate3_562_774 = gate3_620_728 & gate3_647_728;
assign not_304_1107 = ~xor_338_1054;
assign xor_338_1054 = not_480_858 ^ gate3_284_983;
assign gate3_284_983 = gate3_493_774 | gate3_399_857;
assign gate3_399_857 = gate3_569_728 & xor_496_774;
assign xor_496_774 = gate3_563_728 ^ gate3_572_728;
assign gate3_572_728 = lever[11] & lever[32];
assign gate3_563_728 = lever[33] & lever[10];
assign gate3_569_728 = lever[9] & lever[34];
assign gate3_493_774 = gate3_572_728 & gate3_563_728;
assign not_480_858 = ~xor_480_857;
assign xor_480_857 = gate3_659_728 ^ xor_574_774;
assign gate3_334_1054 = not_335_1053 & gate3_284_983;
assign not_335_1053 = ~not_480_858;
assign gate3_261_1233 = xor_315_1108 | not_262_1232;
assign not_262_1232 = ~gate3_216_1182;
assign gate3_179_1453 = gate3_207_1394 & gate3_173_1430;
assign gate3_173_1430 = not_201_1395 | xor_210_1394;
assign xor_210_1394 = gate3_212_1366 ^ not_277_1280;
assign not_277_1280 = ~xor_277_1279;
assign xor_277_1279 = not_270_1234 ^ not_243_1183;
assign gate3_212_1366 = gate3_197_1330 | gate3_241_1279;
assign gate3_241_1279 = gate3_222_1233 & not_242_1278;
assign not_242_1278 = ~xor_286_1108;
assign xor_286_1108 = gate3_527_728 ^ xor_310_1054;
assign gate3_222_1233 = xor_469_774 & not_260_1182;
assign not_260_1182 = ~xor_260_1108;
assign xor_260_1108 = gate3_225_983 ^ xor_280_1054;
assign xor_280_1054 = not_372_858 ^ gate3_228_983;
assign gate3_228_983 = gate3_415_774 | gate3_345_857;
assign gate3_345_857 = gate3_482_728 & xor_418_774;
assign xor_418_774 = gate3_476_728 ^ gate3_485_728;
assign gate3_485_728 = lever[23] & lever[19];
assign gate3_482_728 = lever[25] & lever[17];
assign gate3_415_774 = gate3_470_728 & gate3_488_728;
assign gate3_488_728 = lever[24] & lever[19];
assign gate3_470_728 = lever[18] & lever[23];
assign not_372_858 = ~xor_372_857;
assign xor_372_857 = gate3_515_728 ^ xor_454_774;
assign gate3_225_983 = gate3_436_774 | gate3_357_857;
assign gate3_357_857 = gate3_506_728 & xor_439_774;
assign xor_439_774 = gate3_497_728 ^ gate3_509_728;
assign gate3_509_728 = lever[26] & lever[16];
assign gate3_497_728 = lever[27] & lever[15];
assign gate3_506_728 = lever[28] & lever[14];
assign gate3_436_774 = gate3_497_728 & gate3_509_728;
assign xor_469_774 = gate3_488_728 ^ gate3_524_728;
assign gate3_524_728 = lever[18] & lever[25];
assign gate3_197_1330 = not_244_1280 & not_231_1280;
assign not_231_1280 = ~xor_231_1279;
assign xor_231_1279 = gate3_199_1182 ^ xor_245_1233;
assign xor_245_1233 = xor_279_1108 ^ gate3_202_1182;
assign gate3_202_1182 = gate3_274_1054 | gate3_257_1108;
assign gate3_257_1108 = gate3_225_983 & not_258_1107;
assign not_258_1107 = ~xor_280_1054;
assign gate3_274_1054 = gate3_228_983 & not_275_1053;
assign not_275_1053 = ~not_372_858;
assign xor_279_1108 = not_420_858 ^ xor_301_1054;
assign gate3_199_1182 = gate3_292_1054 & gate3_267_1108;
assign gate3_267_1108 = xor_295_1054 | not_403_858;
assign not_403_858 = ~xor_403_857;
assign xor_403_857 = gate3_569_728 ^ xor_496_774;
assign xor_295_1054 = not_411_858 ^ gate3_234_983;
assign gate3_234_983 = gate3_478_774 | gate3_381_857;
assign gate3_381_857 = gate3_545_728 & xor_484_774;
assign xor_484_774 = gate3_536_728 ^ gate3_548_728;
assign gate3_548_728 = lever[29] & lever[13];
assign gate3_536_728 = lever[30] & lever[12];
assign gate3_545_728 = lever[11] & lever[31];
assign gate3_478_774 = gate3_536_728 & gate3_548_728;
assign not_411_858 = ~xor_411_857;
assign xor_411_857 = gate3_578_728 ^ xor_508_774;
assign gate3_292_1054 = not_411_858 | not_293_1053;
assign not_293_1053 = ~gate3_234_983;
assign not_244_1280 = ~xor_244_1279;
assign xor_244_1279 = gate3_222_1233 ^ xor_286_1108;
assign not_201_1395 = ~xor_201_1394;
assign xor_201_1394 = xor_209_1366 ^ gate3_214_1330;
assign gate3_214_1330 = gate3_255_1233 & not_215_1329;
assign not_215_1329 = ~gate3_253_1279;
assign gate3_253_1279 = not_258_1234 & gate3_656_728;
assign gate3_656_728 = lever[6] & lever[38];
assign not_258_1234 = ~xor_258_1233;
assign xor_258_1233 = gate3_210_1182 ^ xor_306_1108;
assign xor_306_1108 = gate3_278_983 ^ xor_338_1054;
assign gate3_210_1182 = gate3_327_1054 | gate3_294_1108;
assign gate3_294_1108 = gate3_272_983 & not_295_1107;
assign not_295_1107 = ~xor_330_1054;
assign xor_330_1054 = not_465_858 ^ gate3_275_983;
assign gate3_275_983 = gate3_387_857 | gate3_487_774;
assign gate3_487_774 = gate3_557_728 & gate3_560_728;
assign gate3_560_728 = lever[9] & lever[33];
assign gate3_557_728 = lever[10] & lever[32];
assign gate3_387_857 = gate3_554_728 & xor_490_774;
assign xor_490_774 = gate3_557_728 ^ gate3_560_728;
assign gate3_554_728 = lever[8] & lever[34];
assign not_465_858 = ~xor_465_857;
assign xor_465_857 = gate3_644_728 ^ xor_565_774;
assign gate3_272_983 = gate3_535_774 | gate3_441_857;
assign gate3_441_857 = gate3_611_728 & xor_538_774;
assign xor_538_774 = gate3_614_728 ^ gate3_617_728;
assign gate3_617_728 = lever[6] & lever[36];
assign gate3_614_728 = lever[7] & lever[35];
assign gate3_611_728 = lever[5] & lever[37];
assign gate3_535_774 = gate3_614_728 & gate3_617_728;
assign gate3_327_1054 = gate3_275_983 & not_328_1053;
assign not_328_1053 = ~not_465_858;
assign gate3_255_1233 = xor_306_1108 | not_256_1232;
assign not_256_1232 = ~gate3_210_1182;
assign xor_209_1366 = not_266_1280 ^ gate3_217_1330;
assign gate3_217_1330 = gate3_239_1233 | gate3_224_1279;
assign gate3_224_1279 = xor_245_1233 & not_225_1278;
assign not_225_1278 = ~gate3_199_1182;
assign gate3_239_1233 = xor_279_1108 & gate3_202_1182;
assign not_266_1280 = ~xor_266_1279;
assign xor_266_1279 = gate3_668_728 ^ not_264_1234;
assign gate3_207_1394 = not_208_1393 | not_277_1280;
assign not_208_1393 = ~gate3_212_1366;
assign gate3_190_1430 = gate3_205_1366 & gate3_198_1394;
assign gate3_198_1394 = gate3_214_1330 | xor_209_1366;
assign gate3_205_1366 = not_266_1280 | not_206_1365;
assign not_206_1365 = ~gate3_217_1330;
assign gate3_156_1478 = gate3_179_1453 | not_216_1395;
assign not_162_1479 = ~xor_162_1478;
assign xor_162_1478 = gate3_219_1394 ^ xor_183_1453;
assign xor_183_1453 = gate3_193_1430 ^ xor_222_1394;
assign xor_222_1394 = not_231_1367 ^ xor_237_1366;
assign gate3_193_1430 = gate3_213_1394 & gate3_225_1366;
assign gate3_225_1366 = xor_290_1279 | not_226_1365;
assign not_226_1365 = ~gate3_229_1330;
assign gate3_213_1394 = not_219_1367 | xor_228_1366;
assign gate3_219_1394 = gate3_223_1330 & gate3_216_1366;
assign gate3_216_1366 = gate3_220_1330 | xor_226_1330;
assign gate3_223_1330 = not_283_1280 | not_224_1329;
assign not_224_1329 = ~gate3_286_1279;
assign gate3_692_728 = lever[8] & lever[39];
assign gate3_49_1555 = not_162_1479 & not_50_1554;
assign not_50_1554 = ~gate3_157_1528;
assign not_64_1556 = ~xor_64_1555;
assign xor_64_1555 = gate3_65_728 ^ not_76_1529;
assign not_76_1529 = ~xor_76_1528;
assign xor_76_1528 = gate3_42_1503 ^ not_69_1479;
assign not_69_1479 = ~xor_69_1478;
assign xor_69_1478 = gate3_53_1394 ^ xor_85_1453;
assign gate3_42_1503 = gate3_67_1453 & gate3_51_1478;
assign gate3_51_1478 = gate3_219_1394 | not_52_1477;
assign not_52_1477 = ~xor_183_1453;
assign gate3_67_1453 = gate3_193_1430 | xor_222_1394;
assign gate3_65_728 = lever[9] & lever[39];
assign gate3_66_1602 = not_71_1556 & not_67_1601;
assign not_67_1601 = ~gate3_54_1576;
assign gate3_54_1576 = gate3_69_1528 | gate3_56_1555;
assign gate3_56_1555 = gate3_65_728 & not_76_1529;
assign gate3_69_1528 = not_69_1479 & not_70_1527;
assign not_70_1527 = ~gate3_42_1503;
assign not_71_1556 = ~xor_71_1555;
assign xor_71_1555 = gate3_71_728 ^ not_84_1529;
assign gate3_71_1602 = not_72_1601 | not_71_1556;
assign not_72_1601 = ~gate3_54_1576;
assign gate3_1_1885 = gate3_1_1876 | gate3_124_1679;
assign gate3_124_1679 = not_125_1678 | gate3_52_1654;
assign gate3_52_1654 = gate3_84_1628 | gate3_87_1628;
assign gate3_87_1628 = not_64_1556 & not_88_1627;
assign not_88_1627 = ~gate3_57_1602;
assign gate3_84_1628 = not_85_1627 | gate3_66_1602;
assign not_85_1627 = ~gate3_71_1602;
assign not_125_1678 = ~gate3_77_1628;
assign gate3_1_1876 = gate3_62_1628 | gate3_1_1866;
assign gate3_1_1866 = gate3_1_1857 & gate3_59_1693;
assign gate3_59_1693 = gate3_111_1679 & gate3_59_1628;
assign gate3_59_1628 = not_43_1577 | not_60_1627;
assign not_60_1627 = ~gate3_54_1602;
assign gate3_54_1602 = gate3_117_1576 | gate3_133_1555;
assign gate3_133_1555 = not_134_1504 & not_134_1554;
assign not_134_1554 = ~gate3_154_1528;
assign gate3_154_1528 = gate3_147_1478 & gate3_125_1503;
assign gate3_125_1503 = gate3_187_1430 | not_126_1502;
assign not_126_1502 = ~xor_150_1478;
assign xor_150_1478 = not_181_1431 ^ gate3_173_1453;
assign gate3_173_1453 = gate3_185_1394 & gate3_170_1430;
assign gate3_170_1430 = not_191_1395 | xor_195_1394;
assign xor_195_1394 = gate3_190_1366 ^ not_200_1331;
assign not_200_1331 = ~xor_200_1330;
assign xor_200_1330 = not_231_1280 ^ not_244_1280;
assign gate3_190_1366 = gate3_212_1279 | gate3_194_1330;
assign gate3_194_1330 = not_221_1280 & not_218_1280;
assign not_218_1280 = ~xor_218_1279;
assign xor_218_1279 = not_231_1234 ^ gate3_191_1182;
assign gate3_191_1182 = gate3_284_1054 & gate3_264_1108;
assign gate3_264_1108 = not_396_858 | xor_287_1054;
assign xor_287_1054 = gate3_231_983 ^ not_384_858;
assign not_384_858 = ~xor_384_857;
assign xor_384_857 = xor_484_774 ^ gate3_545_728;
assign gate3_231_983 = gate3_472_774 | gate3_378_857;
assign gate3_378_857 = gate3_542_728 & xor_475_774;
assign xor_475_774 = gate3_530_728 ^ gate3_533_728;
assign gate3_533_728 = lever[30] & lever[11];
assign gate3_530_728 = lever[29] & lever[12];
assign gate3_542_728 = lever[10] & lever[31];
assign gate3_472_774 = gate3_530_728 & gate3_533_728;
assign not_396_858 = ~xor_396_857;
assign xor_396_857 = gate3_554_728 ^ xor_490_774;
assign gate3_284_1054 = not_384_858 | not_285_1053;
assign not_285_1053 = ~gate3_231_983;
assign not_231_1234 = ~xor_231_1233;
assign xor_231_1233 = xor_270_1108 ^ gate3_196_1182;
assign gate3_196_1182 = gate3_262_1054 & gate3_248_1108;
assign gate3_248_1108 = xor_265_1054 | not_249_1107;
assign not_249_1107 = ~gate3_216_983;
assign gate3_216_983 = gate3_427_774 | gate3_354_857;
assign gate3_354_857 = gate3_503_728 & xor_430_774;
assign xor_430_774 = gate3_491_728 ^ gate3_494_728;
assign gate3_494_728 = lever[27] & lever[14];
assign gate3_491_728 = lever[26] & lever[15];
assign gate3_503_728 = lever[28] & lever[13];
assign gate3_427_774 = gate3_491_728 & gate3_494_728;
assign xor_265_1054 = not_363_858 ^ gate3_219_983;
assign gate3_219_983 = gate3_406_774 | gate3_336_857;
assign gate3_336_857 = gate3_467_728 & xor_409_774;
assign xor_409_774 = gate3_470_728 ^ gate3_473_728;
assign gate3_473_728 = lever[24] & lever[17];
assign gate3_467_728 = lever[25] & lever[16];
assign gate3_406_774 = gate3_476_728 & gate3_479_728;
assign gate3_479_728 = lever[17] & lever[23];
assign not_363_858 = ~xor_363_857;
assign xor_363_857 = gate3_506_728 ^ xor_439_774;
assign gate3_262_1054 = not_363_858 | not_263_1053;
assign not_263_1053 = ~gate3_219_983;
assign xor_270_1108 = not_403_858 ^ xor_295_1054;
assign not_221_1280 = ~xor_221_1279;
assign xor_221_1279 = gate3_219_1233 ^ not_188_1183;
assign not_188_1183 = ~xor_188_1182;
assign xor_188_1182 = xor_260_1108 ^ xor_469_774;
assign gate3_219_1233 = gate3_245_1108 & gate3_185_1182;
assign gate3_185_1182 = xor_251_1108 | not_186_1181;
assign not_186_1181 = ~xor_254_1108;
assign xor_254_1108 = not_348_858 ^ gate3_259_1054;
assign gate3_259_1054 = gate3_330_857 & gate3_213_983;
assign gate3_213_983 = gate3_394_774 | not_342_858;
assign not_342_858 = ~xor_342_857;
assign xor_342_857 = xor_409_774 ^ gate3_467_728;
assign gate3_394_774 = gate3_461_728 | not_395_773;
assign not_395_773 = ~gate3_464_728;
assign gate3_464_728 = lever[22] & lever[19];
assign gate3_461_728 = lever[21] & lever[18];
assign gate3_330_857 = not_461_774 | not_331_856;
assign not_331_856 = ~gate3_464_728;
assign not_461_774 = ~gate3_461_728;
assign not_348_858 = ~xor_348_857;
assign xor_348_857 = gate3_482_728 ^ xor_418_774;
assign xor_251_1108 = gate3_216_983 ^ xor_265_1054;
assign gate3_245_1108 = gate3_259_1054 | not_348_858;
assign gate3_212_1279 = not_188_1183 & not_213_1278;
assign not_213_1278 = ~gate3_219_1233;
assign not_191_1395 = ~xor_191_1394;
assign xor_191_1394 = gate3_203_1330 ^ xor_196_1366;
assign xor_196_1366 = not_257_1280 ^ gate3_209_1330;
assign gate3_209_1330 = gate3_227_1233 | gate3_215_1279;
assign gate3_215_1279 = not_231_1234 & not_216_1278;
assign not_216_1278 = ~gate3_191_1182;
assign gate3_227_1233 = xor_270_1108 & not_228_1232;
assign not_228_1232 = ~gate3_196_1182;
assign not_257_1280 = ~xor_257_1279;
assign xor_257_1279 = gate3_656_728 ^ not_258_1234;
assign gate3_203_1330 = gate3_248_1233 & not_204_1329;
assign not_204_1329 = ~gate3_250_1279;
assign gate3_250_1279 = gate3_653_728 & not_251_1234;
assign not_251_1234 = ~xor_251_1233;
assign xor_251_1233 = gate3_207_1182 ^ xor_300_1108;
assign xor_300_1108 = gate3_272_983 ^ xor_330_1054;
assign gate3_207_1182 = gate3_313_1054 | gate3_289_1108;
assign gate3_289_1108 = gate3_267_983 & not_290_1107;
assign not_290_1107 = ~xor_324_1054;
assign xor_324_1054 = not_448_858 ^ gate3_261_983;
assign gate3_261_983 = gate3_547_774 | gate3_453_857;
assign gate3_453_857 = gate3_632_728 & xor_550_774;
assign xor_550_774 = gate3_566_728 ^ gate3_626_728;
assign gate3_626_728 = lever[8] & lever[33];
assign gate3_566_728 = lever[32] & lever[9];
assign gate3_632_728 = lever[7] & lever[34];
assign gate3_547_774 = gate3_566_728 & gate3_626_728;
assign not_448_858 = ~xor_448_857;
assign xor_448_857 = gate3_611_728 ^ xor_538_774;
assign gate3_267_983 = gate3_556_774 | gate3_459_857;
assign gate3_459_857 = gate3_641_728 & xor_559_774;
assign xor_559_774 = gate3_623_728 ^ gate3_635_728;
assign gate3_635_728 = lever[36] & lever[5];
assign gate3_623_728 = lever[35] & lever[6];
assign gate3_641_728 = lever[4] & lever[37];
assign gate3_556_774 = gate3_623_728 & gate3_635_728;
assign gate3_313_1054 = gate3_261_983 & not_314_1053;
assign not_314_1053 = ~not_448_858;
assign gate3_653_728 = lever[5] & lever[38];
assign gate3_248_1233 = xor_300_1108 | not_249_1232;
assign not_249_1232 = ~gate3_207_1182;
assign gate3_185_1394 = not_200_1331 | not_186_1393;
assign not_186_1393 = ~gate3_190_1366;
assign not_181_1431 = ~xor_181_1430;
assign xor_181_1430 = not_201_1395 ^ xor_210_1394;
assign gate3_187_1430 = gate3_193_1366 & gate3_188_1394;
assign gate3_188_1394 = gate3_203_1330 | xor_196_1366;
assign gate3_193_1366 = not_257_1280 | not_194_1365;
assign not_194_1365 = ~gate3_209_1330;
assign gate3_147_1478 = gate3_173_1453 | not_181_1431;
assign not_134_1504 = ~xor_134_1503;
assign xor_134_1503 = gate3_190_1430 ^ xor_159_1478;
assign gate3_117_1576 = gate3_689_728 & not_138_1556;
assign not_138_1556 = ~xor_138_1555;
assign xor_138_1555 = gate3_154_1528 ^ not_134_1504;
assign gate3_689_728 = lever[7] & lever[39];
assign not_43_1577 = ~xor_43_1576;
assign xor_43_1576 = not_142_1556 ^ gate3_692_728;
assign gate3_111_1679 = not_127_1577 | not_112_1678;
assign not_112_1678 = ~gate3_132_1654;
assign gate3_132_1654 = gate3_138_1602 | gate3_143_1628;
assign gate3_143_1628 = gate3_62_728 & not_48_1603;
assign not_48_1603 = ~xor_48_1602;
assign xor_48_1602 = gate3_120_1576 ^ not_140_1504;
assign not_140_1504 = ~xor_140_1503;
assign xor_140_1503 = gate3_187_1430 ^ xor_150_1478;
assign gate3_120_1576 = gate3_160_1528 & gate3_147_1555;
assign gate3_147_1555 = gate3_49_1430 | not_148_1554;
assign not_148_1554 = ~xor_57_1528;
assign xor_57_1528 = gate3_137_1503 ^ not_199_1431;
assign not_199_1431 = ~xor_199_1430;
assign xor_199_1430 = not_191_1395 ^ xor_195_1394;
assign gate3_137_1503 = gate3_165_1478 & gate3_192_1453;
assign gate3_192_1453 = not_249_1331 | not_193_1452;
assign not_193_1452 = ~gate3_196_1430;
assign gate3_196_1430 = gate3_227_1394 | gate3_240_1366;
assign gate3_240_1366 = not_275_1183 & not_241_1365;
assign not_241_1365 = ~gate3_246_1330;
assign gate3_246_1330 = gate3_299_1233 & gate3_307_1279;
assign gate3_307_1279 = xor_372_1108 | not_308_1278;
assign not_308_1278 = ~xor_302_1233;
assign xor_302_1233 = not_332_984 ^ gate3_272_1182;
assign gate3_272_1182 = gate3_357_1108 & gate3_385_1054;
assign gate3_385_1054 = not_628_775 | not_386_1053;
assign not_386_1053 = ~gate3_327_983;
assign gate3_327_983 = gate3_537_857 | gate3_622_774;
assign gate3_622_774 = gate3_701_728 & gate3_455_728;
assign gate3_455_728 = lever[21] & lever[19];
assign gate3_701_728 = lever[18] & lever[20];
assign gate3_537_857 = gate3_704_728 & xor_625_774;
assign xor_625_774 = gate3_698_728 ^ gate3_461_728;
assign gate3_698_728 = lever[19] & lever[20];
assign gate3_704_728 = lever[22] & lever[17];
assign not_628_775 = ~xor_628_774;
assign xor_628_774 = gate3_455_728 ^ gate3_458_728;
assign gate3_458_728 = lever[22] & lever[18];
assign gate3_357_1108 = not_543_858 | xor_388_1054;
assign xor_388_1054 = not_628_775 ^ gate3_327_983;
assign not_543_858 = ~xor_543_857;
assign xor_543_857 = gate3_707_728 ^ xor_637_774;
assign xor_637_774 = gate3_479_728 ^ gate3_710_728;
assign gate3_710_728 = lever[24] & lever[16];
assign gate3_707_728 = lever[25] & lever[15];
assign not_332_984 = ~xor_332_983;
assign xor_332_983 = gate3_394_774 ^ not_342_858;
assign xor_372_1108 = gate3_336_983 ^ xor_405_1054;
assign xor_405_1054 = not_552_858 ^ gate3_339_983;
assign gate3_339_983 = gate3_634_774 | gate3_540_857;
assign gate3_540_857 = xor_637_774 & gate3_707_728;
assign gate3_634_774 = gate3_479_728 & gate3_710_728;
assign not_552_858 = ~xor_552_857;
assign xor_552_857 = gate3_503_728 ^ xor_430_774;
assign gate3_336_983 = gate3_646_774 | gate3_549_857;
assign gate3_549_857 = xor_649_774 & gate3_722_728;
assign gate3_722_728 = lever[28] & lever[12];
assign xor_649_774 = gate3_716_728 ^ gate3_500_728;
assign gate3_500_728 = lever[26] & lever[14];
assign gate3_716_728 = lever[13] & lever[27];
assign gate3_646_774 = gate3_500_728 & gate3_716_728;
assign gate3_299_1233 = gate3_272_1182 | not_332_984;
assign not_275_1183 = ~xor_275_1182;
assign xor_275_1182 = xor_251_1108 ^ xor_254_1108;
assign gate3_227_1394 = not_315_1280 & not_243_1367;
assign not_243_1367 = ~xor_243_1366;
assign xor_243_1366 = not_275_1183 ^ gate3_246_1330;
assign not_315_1280 = ~xor_315_1279;
assign xor_315_1279 = gate3_281_1182 ^ xor_310_1233;
assign xor_310_1233 = xor_387_1108 ^ gate3_284_1182;
assign gate3_284_1182 = gate3_398_1054 | gate3_366_1108;
assign gate3_366_1108 = gate3_336_983 & not_367_1107;
assign not_367_1107 = ~xor_405_1054;
assign gate3_398_1054 = gate3_339_983 & not_399_1053;
assign not_399_1053 = ~not_552_858;
assign xor_387_1108 = not_396_858 ^ xor_287_1054;
assign gate3_281_1182 = gate3_410_1054 & gate3_378_1108;
assign gate3_378_1108 = not_567_858 | xor_415_1054;
assign xor_415_1054 = not_564_858 ^ gate3_342_983;
assign gate3_342_983 = gate3_661_774 | gate3_558_857;
assign gate3_558_857 = gate3_731_728 & xor_664_774;
assign xor_664_774 = gate3_539_728 ^ gate3_725_728;
assign gate3_725_728 = lever[30] & lever[10];
assign gate3_539_728 = lever[11] & lever[29];
assign gate3_731_728 = lever[9] & lever[31];
assign gate3_661_774 = gate3_539_728 & gate3_725_728;
assign not_564_858 = ~xor_564_857;
assign xor_564_857 = gate3_542_728 ^ xor_475_774;
assign not_567_858 = ~xor_567_857;
assign xor_567_857 = xor_550_774 ^ gate3_632_728;
assign gate3_410_1054 = not_564_858 | not_411_1053;
assign not_411_1053 = ~gate3_342_983;
assign not_249_1331 = ~xor_249_1330;
assign xor_249_1330 = not_218_1280 ^ not_221_1280;
assign gate3_165_1478 = xor_195_1453 | not_233_1395;
assign not_233_1395 = ~xor_233_1394;
assign xor_233_1394 = gate3_252_1330 ^ xor_254_1366;
assign xor_254_1366 = not_324_1280 ^ gate3_255_1330;
assign gate3_255_1330 = gate3_305_1233 | gate3_310_1279;
assign gate3_310_1279 = xor_310_1233 & not_311_1278;
assign not_311_1278 = ~gate3_281_1182;
assign gate3_305_1233 = xor_387_1108 & gate3_284_1182;
assign not_324_1280 = ~xor_324_1279;
assign xor_324_1279 = gate3_653_728 ^ not_251_1234;
assign gate3_252_1330 = gate3_313_1233 & not_253_1329;
assign not_253_1329 = ~gate3_318_1279;
assign gate3_318_1279 = not_316_1234 & gate3_752_728;
assign gate3_752_728 = lever[4] & lever[38];
assign not_316_1234 = ~xor_316_1233;
assign xor_316_1233 = gate3_288_1182 ^ xor_396_1108;
assign xor_396_1108 = gate3_267_983 ^ xor_324_1054;
assign gate3_288_1182 = gate3_418_1054 | gate3_393_1108;
assign gate3_393_1108 = not_394_1107 & gate3_350_983;
assign gate3_350_983 = gate3_700_774 | gate3_582_857;
assign gate3_582_857 = gate3_749_728 & xor_709_774;
assign xor_709_774 = gate3_638_728 ^ gate3_743_728;
assign gate3_743_728 = lever[4] & lever[36];
assign gate3_638_728 = lever[35] & lever[5];
assign gate3_749_728 = lever[37] & lever[3];
assign gate3_700_774 = gate3_638_728 & gate3_743_728;
assign not_394_1107 = ~xor_426_1054;
assign xor_426_1054 = not_573_858 ^ gate3_345_983;
assign gate3_345_983 = gate3_682_774 | gate3_576_857;
assign gate3_576_857 = gate3_740_728 & xor_697_774;
assign xor_697_774 = gate3_629_728 ^ gate3_734_728;
assign gate3_734_728 = lever[33] & lever[7];
assign gate3_629_728 = lever[8] & lever[32];
assign gate3_740_728 = lever[6] & lever[34];
assign gate3_682_774 = gate3_629_728 & gate3_734_728;
assign not_573_858 = ~xor_573_857;
assign xor_573_857 = gate3_641_728 ^ xor_559_774;
assign gate3_418_1054 = gate3_345_983 & not_419_1053;
assign not_419_1053 = ~not_573_858;
assign gate3_313_1233 = xor_396_1108 | not_314_1232;
assign not_314_1232 = ~gate3_288_1182;
assign xor_195_1453 = gate3_196_1430 ^ not_249_1331;
assign gate3_49_1430 = gate3_246_1366 & gate3_230_1394;
assign gate3_230_1394 = gate3_252_1330 | xor_254_1366;
assign gate3_246_1366 = not_324_1280 | not_247_1365;
assign not_247_1365 = ~gate3_255_1330;
assign gate3_160_1528 = gate3_137_1503 | not_199_1431;
assign gate3_62_728 = lever[6] & lever[39];
assign gate3_138_1602 = not_140_1504 & not_139_1601;
assign not_139_1601 = ~gate3_120_1576;
assign not_127_1577 = ~xor_127_1576;
assign xor_127_1576 = gate3_689_728 ^ not_138_1556;
assign gate3_1_1857 = gate3_1_1849 | xor_108_1679;
assign xor_108_1679 = gate3_132_1654 ^ not_127_1577;
assign gate3_1_1849 = gate3_1_1841 & gate3_45_1706;
assign gate3_45_1706 = gate3_77_1679 & gate3_45_1693;
assign gate3_45_1693 = xor_86_1679 | gate3_94_1679;
assign gate3_94_1679 = not_56_1629 | not_95_1678;
assign not_95_1678 = ~gate3_49_1654;
assign gate3_49_1654 = gate3_51_1602 | gate3_53_1628;
assign gate3_53_1628 = gate3_929_728 & not_147_1603;
assign not_147_1603 = ~xor_147_1602;
assign xor_147_1602 = not_162_1556 ^ gate3_138_1576;
assign gate3_138_1576 = gate3_170_1528 & gate3_153_1555;
assign gate3_153_1555 = gate3_212_1430 | not_154_1554;
assign not_154_1554 = ~xor_173_1528;
assign xor_173_1528 = not_184_1479 ^ gate3_149_1503;
assign gate3_149_1503 = gate3_207_1453 & gate3_175_1478;
assign gate3_175_1478 = not_268_1395 | xor_214_1453;
assign xor_214_1453 = gate3_205_1430 ^ not_275_1395;
assign not_275_1395 = ~xor_275_1394;
assign xor_275_1394 = not_401_1280 ^ xor_293_1366;
assign xor_293_1366 = gate3_285_1330 ^ not_404_1280;
assign not_404_1280 = ~xor_404_1279;
assign xor_404_1279 = xor_302_1233 ^ xor_372_1108;
assign gate3_285_1330 = gate3_349_1233 | not_286_1329;
assign not_286_1329 = ~gate3_360_1279;
assign gate3_360_1279 = not_361_1278 | xor_471_1108;
assign xor_471_1108 = gate3_393_983 ^ xor_491_1054;
assign xor_491_1054 = not_723_858 ^ gate3_398_983;
assign gate3_398_983 = gate3_784_774 | gate3_658_857;
assign gate3_658_857 = gate3_833_728 & xor_787_774;
assign xor_787_774 = gate3_713_728 ^ gate3_800_728;
assign gate3_800_728 = lever[15] & lever[24];
assign gate3_713_728 = lever[23] & lever[16];
assign gate3_833_728 = lever[25] & lever[14];
assign gate3_784_774 = gate3_713_728 & gate3_800_728;
assign not_723_858 = ~xor_723_857;
assign xor_723_857 = gate3_722_728 ^ xor_649_774;
assign gate3_393_983 = gate3_775_774 | gate3_648_857;
assign gate3_648_857 = gate3_830_728 & xor_781_774;
assign xor_781_774 = gate3_719_728 ^ gate3_827_728;
assign gate3_827_728 = lever[27] & lever[12];
assign gate3_719_728 = lever[13] & lever[26];
assign gate3_830_728 = lever[28] & lever[11];
assign gate3_775_774 = gate3_719_728 & gate3_827_728;
assign not_361_1278 = ~not_352_1234;
assign not_352_1234 = ~xor_352_1233;
assign xor_352_1233 = gate3_317_1182 ^ xor_474_1108;
assign xor_474_1108 = not_543_858 ^ xor_388_1054;
assign gate3_317_1182 = gate3_461_1054 & gate3_431_1108;
assign gate3_431_1108 = not_663_858 | xor_464_1054;
assign xor_464_1054 = gate3_377_983 ^ not_666_858;
assign not_666_858 = ~xor_666_857;
assign xor_666_857 = gate3_704_728 ^ xor_625_774;
assign gate3_377_983 = gate3_745_774 | gate3_624_857;
assign gate3_624_857 = gate3_803_728 & xor_754_774;
assign xor_754_774 = gate3_701_728 ^ gate3_776_728;
assign gate3_776_728 = lever[17] & lever[21];
assign gate3_803_728 = lever[22] & lever[16];
assign gate3_745_774 = gate3_461_728 & gate3_773_728;
assign gate3_773_728 = lever[20] & lever[17];
assign not_663_858 = ~xor_663_857;
assign xor_663_857 = gate3_833_728 ^ xor_787_774;
assign gate3_461_1054 = not_666_858 | not_462_1053;
assign not_462_1053 = ~gate3_377_983;
assign gate3_349_1233 = not_350_1232 & xor_474_1108;
assign not_350_1232 = ~gate3_317_1182;
assign not_401_1280 = ~xor_401_1279;
assign xor_401_1279 = gate3_334_1182 ^ xor_393_1233;
assign xor_393_1233 = gate3_338_1182 ^ xor_505_1108;
assign xor_505_1108 = not_567_858 ^ xor_415_1054;
assign gate3_338_1182 = gate3_488_1054 | gate3_463_1108;
assign gate3_463_1108 = gate3_393_983 & not_464_1107;
assign not_464_1107 = ~xor_491_1054;
assign gate3_488_1054 = gate3_398_983 & not_489_1053;
assign not_489_1053 = ~not_723_858;
assign gate3_334_1182 = gate3_482_1054 & gate3_456_1108;
assign gate3_456_1108 = not_714_858 | xor_485_1054;
assign xor_485_1054 = not_720_858 ^ gate3_389_983;
assign gate3_389_983 = gate3_826_774 | gate3_705_857;
assign gate3_705_857 = xor_835_774 & gate3_878_728;
assign gate3_878_728 = lever[8] & lever[31];
assign xor_835_774 = gate3_857_728 ^ gate3_728_728;
assign gate3_728_728 = lever[10] & lever[29];
assign gate3_857_728 = lever[30] & lever[9];
assign gate3_826_774 = gate3_725_728 & gate3_854_728;
assign gate3_854_728 = lever[9] & lever[29];
assign not_720_858 = ~xor_720_857;
assign xor_720_857 = gate3_731_728 ^ xor_664_774;
assign not_714_858 = ~xor_714_857;
assign xor_714_857 = gate3_740_728 ^ xor_697_774;
assign gate3_482_1054 = not_483_1053 | not_720_858;
assign not_483_1053 = ~gate3_389_983;
assign gate3_205_1430 = gate3_263_1366 | gate3_242_1394;
assign gate3_242_1394 = not_357_1280 & xor_266_1366;
assign xor_266_1366 = gate3_262_1330 ^ not_367_1280;
assign not_367_1280 = ~xor_367_1279;
assign xor_367_1279 = xor_471_1108 ^ not_352_1234;
assign gate3_262_1330 = gate3_328_1233 | not_263_1329;
assign not_263_1329 = ~gate3_333_1279;
assign gate3_333_1279 = xor_427_1108 | not_334_1278;
assign not_334_1278 = ~not_331_1234;
assign not_331_1234 = ~xor_331_1233;
assign xor_331_1233 = xor_434_1108 ^ gate3_294_1182;
assign gate3_294_1182 = gate3_436_1054 & gate3_406_1108;
assign gate3_406_1108 = not_612_858 | xor_439_1054;
assign xor_439_1054 = gate3_356_983 ^ not_630_858;
assign not_630_858 = ~xor_630_857;
assign xor_630_857 = gate3_803_728 ^ xor_754_774;
assign gate3_356_983 = gate3_718_774 | gate3_591_857;
assign gate3_591_857 = gate3_770_728 & xor_724_774;
assign xor_724_774 = gate3_761_728 ^ gate3_773_728;
assign gate3_761_728 = lever[16] & lever[21];
assign gate3_770_728 = lever[22] & lever[15];
assign gate3_718_774 = gate3_761_728 & gate3_773_728;
assign not_612_858 = ~xor_612_857;
assign xor_612_857 = gate3_794_728 ^ xor_742_774;
assign xor_742_774 = gate3_788_728 ^ gate3_797_728;
assign gate3_797_728 = lever[23] & lever[15];
assign gate3_788_728 = lever[14] & lever[24];
assign gate3_794_728 = lever[25] & lever[13];
assign gate3_436_1054 = not_630_858 | not_437_1053;
assign not_437_1053 = ~gate3_356_983;
assign xor_434_1108 = not_663_858 ^ xor_464_1054;
assign xor_427_1108 = gate3_368_983 ^ xor_458_1054;
assign xor_458_1054 = not_651_858 ^ gate3_374_983;
assign gate3_374_983 = gate3_736_774 | gate3_609_857;
assign gate3_609_857 = xor_742_774 & gate3_794_728;
assign gate3_736_774 = gate3_788_728 & gate3_797_728;
assign not_651_858 = ~xor_651_857;
assign xor_651_857 = gate3_830_728 ^ xor_781_774;
assign gate3_368_983 = gate3_763_774 | gate3_639_857;
assign gate3_639_857 = gate3_821_728 & xor_772_774;
assign xor_772_774 = gate3_824_728 ^ gate3_812_728;
assign gate3_812_728 = lever[27] & lever[11];
assign gate3_824_728 = lever[26] & lever[12];
assign gate3_821_728 = lever[28] & lever[10];
assign gate3_763_774 = gate3_812_728 & gate3_824_728;
assign gate3_328_1233 = xor_434_1108 & not_329_1232;
assign not_329_1232 = ~gate3_294_1182;
assign not_357_1280 = ~xor_357_1279;
assign xor_357_1279 = gate3_308_1182 ^ xor_346_1233;
assign xor_346_1233 = xor_459_1108 ^ gate3_311_1182;
assign gate3_311_1182 = gate3_454_1054 | gate3_424_1108;
assign gate3_424_1108 = not_425_1107 & gate3_368_983;
assign not_425_1107 = ~xor_458_1054;
assign gate3_454_1054 = gate3_374_983 & not_455_1053;
assign not_455_1053 = ~not_651_858;
assign xor_459_1108 = not_714_858 ^ xor_485_1054;
assign gate3_308_1182 = gate3_476_1054 & gate3_441_1108;
assign gate3_441_1108 = not_702_858 | xor_479_1054;
assign xor_479_1054 = gate3_386_983 ^ not_708_858;
assign not_708_858 = ~xor_708_857;
assign xor_708_857 = gate3_878_728 ^ xor_835_774;
assign gate3_386_983 = gate3_799_774 | gate3_673_857;
assign gate3_673_857 = gate3_851_728 & xor_805_774;
assign xor_805_774 = gate3_842_728 ^ gate3_854_728;
assign gate3_842_728 = lever[30] & lever[8];
assign gate3_851_728 = lever[7] & lever[31];
assign gate3_799_774 = gate3_842_728 & gate3_854_728;
assign not_702_858 = ~xor_702_857;
assign xor_702_857 = gate3_875_728 ^ xor_823_774;
assign xor_823_774 = gate3_737_728 ^ gate3_869_728;
assign gate3_869_728 = lever[6] & lever[33];
assign gate3_737_728 = lever[32] & lever[7];
assign gate3_875_728 = lever[5] & lever[34];
assign gate3_476_1054 = not_708_858 | not_477_1053;
assign not_477_1053 = ~gate3_386_983;
assign gate3_263_1366 = gate3_262_1330 & not_367_1280;
assign not_268_1395 = ~xor_268_1394;
assign xor_268_1394 = gate3_279_1330 ^ xor_284_1366;
assign xor_284_1366 = not_393_1280 ^ gate3_282_1330;
assign gate3_282_1330 = gate3_342_1233 | gate3_351_1279;
assign gate3_351_1279 = xor_346_1233 & not_352_1278;
assign not_352_1278 = ~gate3_308_1182;
assign gate3_342_1233 = xor_459_1108 & gate3_311_1182;
assign not_393_1280 = ~xor_393_1279;
assign xor_393_1279 = gate3_923_728 ^ not_386_1234;
assign not_386_1234 = ~xor_386_1233;
assign xor_386_1233 = gate3_328_1182 ^ xor_501_1108;
assign xor_501_1108 = gate3_350_983 ^ xor_426_1054;
assign gate3_328_1182 = gate3_509_1054 | gate3_493_1108;
assign gate3_493_1108 = gate3_424_983 & not_494_1107;
assign not_494_1107 = ~xor_514_1054;
assign xor_514_1054 = not_754_858 ^ gate3_427_983;
assign gate3_427_983 = gate3_814_774 | gate3_697_857;
assign gate3_697_857 = xor_823_774 & gate3_875_728;
assign gate3_814_774 = gate3_737_728 & gate3_869_728;
assign not_754_858 = ~xor_754_857;
assign xor_754_857 = gate3_749_728 ^ xor_709_774;
assign gate3_424_983 = gate3_865_774 | gate3_747_857;
assign gate3_747_857 = xor_868_774 & gate3_914_728;
assign gate3_914_728 = lever[2] & lever[37];
assign xor_868_774 = gate3_746_728 ^ gate3_893_728;
assign gate3_893_728 = lever[3] & lever[36];
assign gate3_746_728 = lever[4] & lever[35];
assign gate3_865_774 = gate3_893_728 & gate3_746_728;
assign gate3_509_1054 = gate3_427_983 & not_510_1053;
assign not_510_1053 = ~not_754_858;
assign gate3_923_728 = lever[38] & lever[3];
assign gate3_279_1330 = gate3_365_1233 & not_280_1329;
assign not_280_1329 = ~gate3_373_1279;
assign gate3_373_1279 = not_374_1234 & gate3_920_728;
assign gate3_920_728 = lever[2] & lever[38];
assign not_374_1234 = ~xor_374_1233;
assign xor_374_1233 = xor_498_1108 ^ gate3_325_1182;
assign gate3_325_1182 = gate3_484_1108 | gate3_503_1054;
assign gate3_503_1054 = gate3_416_983 & not_504_1053;
assign not_504_1053 = ~not_750_858;
assign not_750_858 = ~xor_750_857;
assign xor_750_857 = gate3_914_728 ^ xor_868_774;
assign gate3_416_983 = gate3_679_857 | gate3_808_774;
assign gate3_808_774 = gate3_863_728 & gate3_866_728;
assign gate3_866_728 = lever[6] & lever[32];
assign gate3_863_728 = lever[33] & lever[5];
assign gate3_679_857 = gate3_860_728 & xor_811_774;
assign xor_811_774 = gate3_863_728 ^ gate3_866_728;
assign gate3_860_728 = lever[4] & lever[34];
assign gate3_484_1108 = not_485_1107 & gate3_413_983;
assign gate3_413_983 = gate3_838_774 | gate3_729_857;
assign gate3_729_857 = gate3_881_728 & xor_841_774;
assign xor_841_774 = gate3_884_728 ^ gate3_887_728;
assign gate3_887_728 = lever[3] & lever[35];
assign gate3_884_728 = lever[2] & lever[36];
assign gate3_881_728 = lever[1] & lever[37];
assign gate3_838_774 = gate3_884_728 & gate3_887_728;
assign not_485_1107 = ~xor_506_1054;
assign xor_506_1054 = not_750_858 ^ gate3_416_983;
assign xor_498_1108 = gate3_424_983 ^ xor_514_1054;
assign gate3_365_1233 = xor_498_1108 | not_366_1232;
assign not_366_1232 = ~gate3_325_1182;
assign gate3_207_1453 = not_275_1395 | not_208_1452;
assign not_208_1452 = ~gate3_205_1430;
assign not_184_1479 = ~xor_184_1478;
assign xor_184_1478 = not_283_1395 ^ xor_224_1453;
assign xor_224_1453 = gate3_224_1430 ^ not_286_1395;
assign not_286_1395 = ~xor_286_1394;
assign xor_286_1394 = not_315_1280 ^ not_243_1367;
assign gate3_224_1430 = gate3_290_1366 | gate3_272_1394;
assign gate3_272_1394 = not_401_1280 & xor_293_1366;
assign gate3_290_1366 = gate3_285_1330 & not_404_1280;
assign not_283_1395 = ~xor_283_1394;
assign xor_283_1394 = gate3_288_1330 ^ xor_300_1366;
assign xor_300_1366 = not_408_1280 ^ gate3_292_1330;
assign gate3_292_1330 = gate3_389_1233 | gate3_398_1279;
assign gate3_398_1279 = xor_393_1233 & not_399_1278;
assign not_399_1278 = ~gate3_334_1182;
assign gate3_389_1233 = gate3_338_1182 & xor_505_1108;
assign not_408_1280 = ~xor_408_1279;
assign xor_408_1279 = gate3_752_728 ^ not_316_1234;
assign gate3_288_1330 = gate3_379_1233 & not_289_1329;
assign not_289_1329 = ~gate3_387_1279;
assign gate3_387_1279 = gate3_923_728 & not_386_1234;
assign gate3_379_1233 = xor_501_1108 | not_380_1232;
assign not_380_1232 = ~gate3_328_1182;
assign gate3_212_1430 = gate3_281_1366 & gate3_265_1394;
assign gate3_265_1394 = gate3_279_1330 | xor_284_1366;
assign gate3_281_1366 = not_393_1280 | not_282_1365;
assign not_282_1365 = ~gate3_282_1330;
assign gate3_170_1528 = gate3_149_1503 | not_184_1479;
assign not_162_1556 = ~xor_162_1555;
assign xor_162_1555 = gate3_227_1430 ^ xor_176_1528;
assign xor_176_1528 = gate3_152_1503 ^ not_194_1479;
assign not_194_1479 = ~xor_194_1478;
assign xor_194_1478 = xor_195_1453 ^ not_233_1395;
assign gate3_152_1503 = gate3_221_1453 & gate3_181_1478;
assign gate3_181_1478 = not_283_1395 | xor_224_1453;
assign gate3_221_1453 = not_286_1395 | not_222_1452;
assign not_222_1452 = ~gate3_224_1430;
assign gate3_227_1430 = gate3_296_1366 & gate3_278_1394;
assign gate3_278_1394 = gate3_288_1330 | xor_300_1366;
assign gate3_296_1366 = not_297_1365 | not_408_1280;
assign not_297_1365 = ~gate3_292_1330;
assign gate3_929_728 = lever[4] & lever[39];
assign gate3_51_1602 = not_162_1556 & not_52_1601;
assign not_52_1601 = ~gate3_138_1576;
assign not_56_1629 = ~xor_56_1628;
assign xor_56_1628 = gate3_59_728 ^ not_45_1603;
assign not_45_1603 = ~xor_45_1602;
assign xor_45_1602 = gate3_40_1576 ^ not_46_1556;
assign not_46_1556 = ~xor_46_1555;
assign xor_46_1555 = gate3_49_1430 ^ xor_57_1528;
assign gate3_40_1576 = gate3_54_1528 & gate3_43_1555;
assign gate3_43_1555 = gate3_227_1430 | not_44_1554;
assign not_44_1554 = ~xor_176_1528;
assign gate3_54_1528 = gate3_152_1503 | not_194_1479;
assign gate3_59_728 = lever[5] & lever[39];
assign xor_86_1679 = gate3_43_1654 ^ not_47_1629;
assign not_47_1629 = ~xor_47_1628;
assign xor_47_1628 = not_48_1603 ^ gate3_62_728;
assign gate3_43_1654 = gate3_39_1602 | gate3_44_1628;
assign gate3_44_1628 = not_45_1603 & gate3_59_728;
assign gate3_39_1602 = not_40_1601 & not_46_1556;
assign not_40_1601 = ~gate3_40_1576;
assign gate3_77_1679 = not_78_1678 | not_47_1629;
assign not_78_1678 = ~gate3_43_1654;
assign gate3_1_1841 = gate3_1_1834 | gate3_32_1714;
assign gate3_32_1714 = xor_86_1679 | gate3_16_1706;
assign gate3_16_1706 = not_94_1693 | gate3_105_1679;
assign gate3_105_1679 = not_56_1629 & not_106_1678;
assign not_106_1678 = ~gate3_49_1654;
assign not_94_1693 = ~gate3_94_1679;
assign gate3_1_1834 = gate3_1_1827 & gate3_71_1679;
assign gate3_71_1679 = not_72_1678 | not_152_1629;
assign not_152_1629 = ~xor_152_1628;
assign xor_152_1628 = gate3_929_728 ^ not_147_1603;
assign not_72_1678 = ~gate3_135_1654;
assign gate3_135_1654 = gate3_141_1602 | gate3_146_1628;
assign gate3_146_1628 = not_144_1603 & gate3_926_728;
assign gate3_926_728 = lever[3] & lever[39];
assign not_144_1603 = ~xor_144_1602;
assign xor_144_1602 = gate3_130_1576 ^ not_156_1556;
assign not_156_1556 = ~xor_156_1555;
assign xor_156_1555 = gate3_212_1430 ^ xor_173_1528;
assign gate3_130_1576 = gate3_164_1528 & gate3_150_1555;
assign gate3_150_1555 = gate3_209_1430 | not_151_1554;
assign not_151_1554 = ~xor_167_1528;
assign xor_167_1528 = gate3_145_1503 ^ not_178_1479;
assign not_178_1479 = ~xor_178_1478;
assign xor_178_1478 = not_268_1395 ^ xor_214_1453;
assign gate3_145_1503 = gate3_201_1453 & gate3_172_1478;
assign gate3_172_1478 = not_259_1395 | xor_204_1453;
assign xor_204_1453 = gate3_202_1430 ^ not_251_1395;
assign not_251_1395 = ~xor_251_1394;
assign xor_251_1394 = not_357_1280 ^ xor_266_1366;
assign gate3_202_1430 = gate3_236_1394 | gate3_257_1366;
assign gate3_257_1366 = gate3_259_1330 & not_338_1280;
assign not_338_1280 = ~xor_338_1279;
assign xor_338_1279 = xor_427_1108 ^ not_331_1234;
assign gate3_259_1330 = gate3_322_1233 | not_260_1329;
assign not_260_1329 = ~gate3_330_1279;
assign gate3_330_1279 = not_331_1278 | xor_420_1108;
assign xor_420_1108 = gate3_359_983 ^ xor_451_1054;
assign xor_451_1054 = not_642_858 ^ gate3_365_983;
assign gate3_365_983 = gate3_727_774 | gate3_600_857;
assign gate3_600_857 = gate3_779_728 & xor_733_774;
assign xor_733_774 = gate3_782_728 ^ gate3_785_728;
assign gate3_785_728 = lever[23] & lever[14];
assign gate3_782_728 = lever[24] & lever[13];
assign gate3_779_728 = lever[25] & lever[12];
assign gate3_727_774 = gate3_782_728 & gate3_785_728;
assign not_642_858 = ~xor_642_857;
assign xor_642_857 = gate3_821_728 ^ xor_772_774;
assign gate3_359_983 = gate3_757_774 | gate3_636_857;
assign gate3_636_857 = xor_760_774 & gate3_818_728;
assign gate3_818_728 = lever[9] & lever[28];
assign xor_760_774 = gate3_806_728 ^ gate3_809_728;
assign gate3_809_728 = lever[26] & lever[11];
assign gate3_806_728 = lever[27] & lever[10];
assign gate3_757_774 = gate3_806_728 & gate3_809_728;
assign not_331_1278 = ~not_325_1234;
assign not_325_1234 = ~xor_325_1233;
assign xor_325_1233 = xor_412_1108 ^ gate3_291_1182;
assign gate3_291_1182 = gate3_429_1054 & gate3_403_1108;
assign gate3_403_1108 = not_603_858 | xor_432_1054;
assign xor_432_1054 = gate3_353_983 ^ not_594_858;
assign not_594_858 = ~xor_594_857;
assign xor_594_857 = gate3_770_728 ^ xor_724_774;
assign gate3_353_983 = gate3_712_774 | gate3_585_857;
assign gate3_585_857 = gate3_767_728 & xor_715_774;
assign xor_715_774 = gate3_755_728 ^ gate3_758_728;
assign gate3_758_728 = lever[20] & lever[16];
assign gate3_755_728 = lever[21] & lever[15];
assign gate3_767_728 = lever[22] & lever[14];
assign gate3_712_774 = gate3_755_728 & gate3_758_728;
assign not_603_858 = ~xor_603_857;
assign xor_603_857 = gate3_779_728 ^ xor_733_774;
assign gate3_429_1054 = not_430_1053 | not_594_858;
assign not_430_1053 = ~gate3_353_983;
assign xor_412_1108 = not_612_858 ^ xor_439_1054;
assign gate3_322_1233 = xor_412_1108 & not_323_1232;
assign not_323_1232 = ~gate3_291_1182;
assign gate3_236_1394 = not_347_1280 & xor_260_1366;
assign xor_260_1366 = gate3_259_1330 ^ not_338_1280;
assign not_347_1280 = ~xor_347_1279;
assign xor_347_1279 = gate3_297_1182 ^ xor_339_1233;
assign xor_339_1233 = xor_450_1108 ^ gate3_302_1182;
assign gate3_302_1182 = gate3_448_1054 | gate3_415_1108;
assign gate3_415_1108 = gate3_359_983 & not_416_1107;
assign not_416_1107 = ~xor_451_1054;
assign gate3_448_1054 = gate3_365_983 & not_449_1053;
assign not_449_1053 = ~not_642_858;
assign xor_450_1108 = not_702_858 ^ xor_479_1054;
assign gate3_297_1182 = gate3_467_1054 & gate3_438_1108;
assign gate3_438_1108 = not_684_858 | xor_471_1054;
assign xor_471_1054 = not_676_858 ^ gate3_380_983;
assign gate3_380_983 = gate3_790_774 | gate3_670_857;
assign gate3_670_857 = gate3_848_728 & xor_796_774;
assign xor_796_774 = gate3_836_728 ^ gate3_839_728;
assign gate3_839_728 = lever[8] & lever[29];
assign gate3_836_728 = lever[30] & lever[7];
assign gate3_848_728 = lever[6] & lever[31];
assign gate3_790_774 = gate3_836_728 & gate3_839_728;
assign not_676_858 = ~xor_676_857;
assign xor_676_857 = gate3_851_728 ^ xor_805_774;
assign not_684_858 = ~xor_684_857;
assign xor_684_857 = gate3_860_728 ^ xor_811_774;
assign gate3_467_1054 = not_676_858 | not_468_1053;
assign not_468_1053 = ~gate3_380_983;
assign not_259_1395 = ~xor_259_1394;
assign xor_259_1394 = gate3_268_1330 ^ xor_273_1366;
assign xor_273_1366 = not_384_1280 ^ gate3_271_1330;
assign gate3_271_1330 = gate3_336_1233 | gate3_344_1279;
assign gate3_344_1279 = not_345_1278 & xor_339_1233;
assign not_345_1278 = ~gate3_297_1182;
assign gate3_336_1233 = xor_450_1108 & gate3_302_1182;
assign not_384_1280 = ~xor_384_1279;
assign xor_384_1279 = gate3_920_728 ^ not_374_1234;
assign gate3_268_1330 = not_269_1329 & gate3_355_1233;
assign gate3_355_1233 = xor_490_1108 | not_356_1232;
assign not_356_1232 = ~gate3_322_1182;
assign gate3_322_1182 = gate3_496_1054 | gate3_478_1108;
assign gate3_478_1108 = gate3_408_983 & not_479_1107;
assign not_479_1107 = ~xor_499_1054;
assign xor_499_1054 = not_732_858 ^ gate3_405_983;
assign gate3_405_983 = gate3_844_774 | gate3_738_857;
assign gate3_738_857 = gate3_902_728 & xor_853_774;
assign xor_853_774 = gate3_872_728 ^ gate3_896_728;
assign gate3_896_728 = lever[33] & lever[4];
assign gate3_872_728 = lever[32] & lever[5];
assign gate3_902_728 = lever[3] & lever[34];
assign gate3_844_774 = gate3_872_728 & gate3_896_728;
assign not_732_858 = ~xor_732_857;
assign xor_732_857 = gate3_881_728 ^ xor_841_774;
assign gate3_408_983 = gate3_856_774 | gate3_741_857;
assign gate3_741_857 = gate3_911_728 & xor_862_774;
assign xor_862_774 = gate3_890_728 ^ gate3_905_728;
assign gate3_905_728 = lever[1] & lever[36];
assign gate3_890_728 = lever[2] & lever[35];
assign gate3_911_728 = lever[37] & lever[0];
assign gate3_856_774 = gate3_890_728 & gate3_905_728;
assign gate3_496_1054 = gate3_405_983 & not_497_1053;
assign not_497_1053 = ~not_732_858;
assign xor_490_1108 = gate3_413_983 ^ xor_506_1054;
assign not_269_1329 = ~gate3_370_1279;
assign gate3_370_1279 = not_359_1234 & gate3_917_728;
assign gate3_917_728 = lever[1] & lever[38];
assign not_359_1234 = ~xor_359_1233;
assign xor_359_1233 = xor_490_1108 ^ gate3_322_1182;
assign gate3_201_1453 = not_202_1452 | not_251_1395;
assign not_202_1452 = ~gate3_202_1430;
assign gate3_209_1430 = gate3_270_1366 & gate3_254_1394;
assign gate3_254_1394 = gate3_268_1330 | xor_273_1366;
assign gate3_270_1366 = not_384_1280 | not_271_1365;
assign not_271_1365 = ~gate3_271_1330;
assign gate3_164_1528 = gate3_145_1503 | not_178_1479;
assign gate3_141_1602 = not_156_1556 & not_142_1601;
assign not_142_1601 = ~gate3_130_1576;
assign gate3_1_1827 = gate3_1_1819 | xor_64_1679;
assign xor_64_1679 = gate3_135_1654 ^ not_152_1629;
assign gate3_1_1819 = gate3_1_1813 & gate3_57_1679;
assign gate3_57_1679 = not_164_1629 | not_58_1678;
assign not_58_1678 = ~gate3_138_1654;
assign gate3_138_1654 = gate3_158_1628 | gate3_150_1602;
assign gate3_150_1602 = not_151_1601 & not_172_1556;
assign not_172_1556 = ~xor_172_1555;
assign xor_172_1555 = gate3_209_1430 ^ xor_167_1528;
assign not_151_1601 = ~gate3_142_1576;
assign gate3_142_1576 = gate3_179_1528 & gate3_166_1555;
assign gate3_166_1555 = gate3_235_1430 | not_167_1554;
assign not_167_1554 = ~xor_182_1528;
assign xor_182_1528 = gate3_158_1503 ^ not_203_1479;
assign not_203_1479 = ~xor_203_1478;
assign xor_203_1478 = xor_204_1453 ^ not_259_1395;
assign gate3_158_1503 = gate3_229_1453 & gate3_197_1478;
assign gate3_197_1478 = xor_305_1394 | xor_237_1453;
assign xor_237_1453 = gate3_230_1430 ^ not_298_1395;
assign not_298_1395 = ~xor_298_1394;
assign xor_298_1394 = not_347_1280 ^ xor_260_1366;
assign gate3_230_1430 = gate3_303_1366 | gate3_292_1394;
assign gate3_292_1394 = not_422_1280 & not_293_1393;
assign not_293_1393 = ~not_306_1367;
assign not_306_1367 = ~xor_306_1366;
assign xor_306_1366 = not_416_1280 ^ gate3_295_1330;
assign gate3_295_1330 = gate3_396_1233 | gate3_411_1279;
assign gate3_411_1279 = not_525_1109 & not_403_1234;
assign not_403_1234 = ~xor_403_1233;
assign xor_403_1233 = gate3_341_1182 ^ xor_514_1108;
assign xor_514_1108 = not_603_858 ^ xor_432_1054;
assign gate3_341_1182 = gate3_517_1054 & gate3_511_1108;
assign gate3_511_1108 = not_771_858 | xor_520_1054;
assign xor_520_1054 = not_765_858 ^ gate3_431_983;
assign gate3_431_983 = gate3_871_774 | gate3_759_857;
assign gate3_759_857 = gate3_938_728 & xor_883_774;
assign xor_883_774 = gate3_764_728 ^ gate3_932_728;
assign gate3_932_728 = lever[21] & lever[14];
assign gate3_764_728 = lever[15] & lever[20];
assign gate3_938_728 = lever[22] & lever[13];
assign gate3_871_774 = gate3_764_728 & gate3_932_728;
assign not_765_858 = ~xor_765_857;
assign xor_765_857 = gate3_767_728 ^ xor_715_774;
assign not_771_858 = ~xor_771_857;
assign xor_771_857 = gate3_941_728 ^ xor_889_774;
assign xor_889_774 = gate3_944_728 ^ gate3_791_728;
assign gate3_791_728 = lever[13] & lever[23];
assign gate3_944_728 = lever[12] & lever[24];
assign gate3_941_728 = lever[25] & lever[11];
assign gate3_517_1054 = not_765_858 | not_518_1053;
assign not_518_1053 = ~gate3_431_983;
assign not_525_1109 = ~xor_525_1108;
assign xor_525_1108 = gate3_434_983 ^ xor_529_1054;
assign xor_529_1054 = gate3_437_983 ^ not_780_858;
assign not_780_858 = ~xor_780_857;
assign xor_780_857 = gate3_818_728 ^ xor_760_774;
assign gate3_437_983 = gate3_886_774 | gate3_768_857;
assign gate3_768_857 = xor_889_774 & gate3_941_728;
assign gate3_886_774 = gate3_791_728 & gate3_944_728;
assign gate3_434_983 = gate3_892_774 | gate3_777_857;
assign gate3_777_857 = gate3_956_728 & xor_895_774;
assign xor_895_774 = gate3_815_728 ^ gate3_950_728;
assign gate3_950_728 = lever[27] & lever[9];
assign gate3_815_728 = lever[26] & lever[10];
assign gate3_956_728 = lever[8] & lever[28];
assign gate3_892_774 = gate3_815_728 & gate3_950_728;
assign gate3_396_1233 = xor_514_1108 & not_397_1232;
assign not_397_1232 = ~gate3_341_1182;
assign not_416_1280 = ~xor_416_1279;
assign xor_416_1279 = xor_420_1108 ^ not_325_1234;
assign not_422_1280 = ~xor_422_1279;
assign xor_422_1279 = gate3_344_1182 ^ not_411_1234;
assign not_411_1234 = ~xor_411_1233;
assign xor_411_1233 = xor_534_1108 ^ gate3_347_1182;
assign gate3_347_1182 = gate3_523_1054 & gate3_519_1108;
assign gate3_519_1108 = not_520_1107 | xor_529_1054;
assign not_520_1107 = ~gate3_434_983;
assign gate3_523_1054 = not_780_858 | not_524_1053;
assign not_524_1053 = ~gate3_437_983;
assign xor_534_1108 = not_684_858 ^ xor_471_1054;
assign gate3_344_1182 = gate3_532_1054 & gate3_528_1108;
assign gate3_528_1108 = not_795_858 | xor_538_1054;
assign xor_538_1054 = gate3_440_983 ^ not_792_858;
assign not_792_858 = ~xor_792_857;
assign xor_792_857 = gate3_848_728 ^ xor_796_774;
assign gate3_440_983 = gate3_898_774 | gate3_786_857;
assign gate3_786_857 = gate3_965_728 & xor_904_774;
assign xor_904_774 = gate3_845_728 ^ gate3_959_728;
assign gate3_959_728 = lever[30] & lever[6];
assign gate3_845_728 = lever[29] & lever[7];
assign gate3_965_728 = lever[5] & lever[31];
assign gate3_898_774 = gate3_845_728 & gate3_959_728;
assign not_795_858 = ~xor_795_857;
assign xor_795_857 = gate3_902_728 ^ xor_853_774;
assign gate3_532_1054 = not_533_1053 | not_792_858;
assign not_533_1053 = ~gate3_440_983;
assign gate3_303_1366 = gate3_295_1330 & not_416_1280;
assign xor_305_1394 = gate3_298_1330 ^ xor_312_1366;
assign xor_312_1366 = not_429_1280 ^ gate3_303_1330;
assign gate3_303_1330 = gate3_406_1233 | gate3_419_1279;
assign gate3_419_1279 = not_411_1234 & not_420_1278;
assign not_420_1278 = ~gate3_344_1182;
assign gate3_406_1233 = not_407_1232 & xor_534_1108;
assign not_407_1232 = ~gate3_347_1182;
assign not_429_1280 = ~xor_429_1279;
assign xor_429_1279 = gate3_917_728 ^ not_359_1234;
assign gate3_298_1330 = gate3_414_1233 | gate3_426_1279;
assign gate3_426_1279 = xor_417_1233 & gate3_983_728;
assign gate3_983_728 = lever[38] & lever[0];
assign xor_417_1233 = not_537_1109 ^ gate3_351_1182;
assign gate3_351_1182 = gate3_541_1054 & gate3_543_1108;
assign gate3_543_1108 = gate3_545_1054 | gate3_934_774;
assign gate3_934_774 = gate3_905_728 & gate3_980_728;
assign gate3_980_728 = lever[35] & lever[0];
assign gate3_545_1054 = gate3_450_983 & not_546_1053;
assign not_546_1053 = ~not_801_858;
assign not_801_858 = ~xor_801_857;
assign xor_801_857 = gate3_911_728 ^ xor_862_774;
assign gate3_450_983 = gate3_907_774 | gate3_804_857;
assign gate3_804_857 = gate3_974_728 & xor_931_774;
assign xor_931_774 = gate3_968_728 ^ gate3_899_728;
assign gate3_899_728 = lever[32] & lever[4];
assign gate3_968_728 = lever[33] & lever[3];
assign gate3_974_728 = lever[2] & lever[34];
assign gate3_907_774 = gate3_899_728 & gate3_968_728;
assign gate3_541_1054 = gate3_450_983 | not_542_1053;
assign not_542_1053 = ~not_801_858;
assign not_537_1109 = ~xor_537_1108;
assign xor_537_1108 = gate3_408_983 ^ xor_499_1054;
assign gate3_414_1233 = gate3_351_1182 & not_537_1109;
assign gate3_229_1453 = not_298_1395 | not_230_1452;
assign not_230_1452 = ~gate3_230_1430;
assign gate3_235_1430 = gate3_309_1366 & gate3_301_1394;
assign gate3_301_1394 = xor_312_1366 | not_302_1393;
assign not_302_1393 = ~gate3_298_1330;
assign gate3_309_1366 = not_429_1280 | not_310_1365;
assign not_310_1365 = ~gate3_303_1330;
assign gate3_179_1528 = gate3_158_1503 | not_203_1479;
assign gate3_158_1628 = gate3_986_728 & not_153_1603;
assign not_153_1603 = ~xor_153_1602;
assign xor_153_1602 = not_172_1556 ^ gate3_142_1576;
assign gate3_986_728 = lever[2] & lever[39];
assign not_164_1629 = ~xor_164_1628;
assign xor_164_1628 = gate3_926_728 ^ not_144_1603;
assign gate3_1_1813 = gate3_1_1805 | xor_54_1679;
assign xor_54_1679 = gate3_138_1654 ^ not_164_1629;
assign gate3_1_1805 = gate3_1_1800 & gate3_4_1706;
assign gate3_4_1706 = gate3_49_1679 & gate3_4_1693;
assign gate3_4_1693 = xor_43_1679 | gate3_46_1679;
assign gate3_46_1679 = not_183_1629 | not_47_1678;
assign not_47_1678 = ~gate3_144_1654;
assign gate3_144_1654 = gate3_180_1628 | gate3_162_1602;
assign gate3_162_1602 = gate3_150_1576 & not_193_1556;
assign not_193_1556 = ~xor_193_1555;
assign xor_193_1555 = gate3_241_1430 ^ not_188_1529;
assign not_188_1529 = ~xor_188_1528;
assign xor_188_1528 = xor_217_1478 ^ gate3_164_1503;
assign gate3_164_1503 = gate3_243_1453 & gate3_214_1478;
assign gate3_214_1478 = xor_249_1453 | not_325_1395;
assign not_325_1395 = ~xor_325_1394;
assign xor_325_1394 = gate3_363_1182 ^ xor_326_1366;
assign xor_326_1366 = gate3_309_1330 ^ not_456_1280;
assign not_456_1280 = ~xor_456_1279;
assign xor_456_1279 = gate3_983_728 ^ xor_417_1233;
assign gate3_309_1330 = gate3_432_1233 | gate3_445_1279;
assign gate3_445_1279 = xor_435_1233 & not_446_1278;
assign not_446_1278 = ~gate3_357_1182;
assign gate3_357_1182 = gate3_565_1054 & gate3_562_1108;
assign gate3_562_1108 = not_846_858 | xor_569_1054;
assign xor_569_1054 = not_840_858 ^ gate3_462_983;
assign gate3_462_983 = gate3_967_774 | gate3_834_857;
assign gate3_834_857 = gate3_1022_728 & xor_970_774;
assign xor_970_774 = gate3_962_728 ^ gate3_1016_728;
assign gate3_1016_728 = lever[30] & lever[5];
assign gate3_962_728 = lever[29] & lever[6];
assign gate3_1022_728 = lever[4] & lever[31];
assign gate3_967_774 = gate3_962_728 & gate3_1016_728;
assign not_840_858 = ~xor_840_857;
assign xor_840_857 = gate3_965_728 ^ xor_904_774;
assign not_846_858 = ~xor_846_857;
assign xor_846_857 = gate3_974_728 ^ xor_931_774;
assign gate3_565_1054 = not_840_858 | not_566_1053;
assign not_566_1053 = ~gate3_462_983;
assign xor_435_1233 = xor_567_1108 ^ gate3_360_1182;
assign gate3_360_1182 = gate3_556_1054 | gate3_553_1108;
assign gate3_553_1108 = gate3_456_983 & not_554_1107;
assign not_554_1107 = ~xor_562_1054;
assign xor_562_1054 = not_831_858 ^ gate3_459_983;
assign gate3_459_983 = gate3_819_857 | gate3_949_774;
assign gate3_949_774 = gate3_947_728 & gate3_1001_728;
assign gate3_1001_728 = lever[24] & lever[11];
assign gate3_947_728 = lever[12] & lever[23];
assign gate3_819_857 = gate3_998_728 & xor_952_774;
assign xor_952_774 = gate3_947_728 ^ gate3_1001_728;
assign gate3_998_728 = lever[25] & lever[10];
assign not_831_858 = ~xor_831_857;
assign xor_831_857 = gate3_956_728 ^ xor_895_774;
assign gate3_456_983 = gate3_958_774 | gate3_828_857;
assign gate3_828_857 = xor_961_774 & gate3_1013_728;
assign gate3_1013_728 = lever[7] & lever[28];
assign xor_961_774 = gate3_1007_728 ^ gate3_953_728;
assign gate3_953_728 = lever[26] & lever[9];
assign gate3_1007_728 = lever[8] & lever[27];
assign gate3_958_774 = gate3_953_728 & gate3_1007_728;
assign gate3_556_1054 = gate3_459_983 & not_557_1053;
assign not_557_1053 = ~not_831_858;
assign xor_567_1108 = not_795_858 ^ xor_538_1054;
assign gate3_432_1233 = xor_567_1108 & gate3_360_1182;
assign gate3_363_1182 = not_572_1108 | xor_575_1054;
assign xor_575_1054 = not_801_858 ^ gate3_450_983;
assign not_572_1108 = ~gate3_572_1054;
assign gate3_572_1054 = xor_976_774 & gate3_467_983;
assign gate3_467_983 = gate3_988_774 | gate3_849_857;
assign gate3_849_857 = xor_991_774 & gate3_1031_728;
assign gate3_1031_728 = lever[34] & lever[1];
assign xor_991_774 = gate3_1025_728 ^ gate3_971_728;
assign gate3_971_728 = lever[3] & lever[32];
assign gate3_1025_728 = lever[2] & lever[33];
assign gate3_988_774 = gate3_971_728 & gate3_1025_728;
assign xor_976_774 = gate3_908_728 ^ gate3_977_728;
assign gate3_977_728 = lever[0] & lever[36];
assign gate3_908_728 = lever[1] & lever[35];
assign xor_249_1453 = xor_314_1394 ^ gate3_238_1430;
assign gate3_238_1430 = gate3_317_1366 | gate3_311_1394;
assign gate3_311_1394 = not_450_1280 & xor_320_1366;
assign xor_320_1366 = xor_440_1279 ^ gate3_306_1330;
assign gate3_306_1330 = gate3_424_1233 | not_307_1329;
assign not_307_1329 = ~gate3_434_1279;
assign gate3_434_1279 = xor_558_1108 | not_435_1278;
assign not_435_1278 = ~not_429_1234;
assign not_429_1234 = ~xor_429_1233;
assign xor_429_1233 = xor_550_1108 ^ gate3_354_1182;
assign gate3_354_1182 = gate3_548_1054 & gate3_546_1108;
assign gate3_546_1108 = not_822_858 | xor_551_1054;
assign xor_551_1054 = gate3_453_983 ^ not_816_858;
assign not_816_858 = ~xor_816_857;
assign xor_816_857 = gate3_938_728 ^ xor_883_774;
assign gate3_453_983 = gate3_943_774 | gate3_810_857;
assign gate3_810_857 = gate3_995_728 & xor_946_774;
assign xor_946_774 = gate3_935_728 ^ gate3_989_728;
assign gate3_989_728 = lever[13] & lever[21];
assign gate3_935_728 = lever[20] & lever[14];
assign gate3_995_728 = lever[22] & lever[12];
assign gate3_943_774 = gate3_935_728 & gate3_989_728;
assign not_822_858 = ~xor_822_857;
assign xor_822_857 = gate3_998_728 ^ xor_952_774;
assign gate3_548_1054 = not_816_858 | not_549_1053;
assign not_549_1053 = ~gate3_453_983;
assign xor_550_1108 = not_771_858 ^ xor_520_1054;
assign xor_558_1108 = gate3_456_983 ^ xor_562_1054;
assign gate3_424_1233 = xor_550_1108 & not_425_1232;
assign not_425_1232 = ~gate3_354_1182;
assign xor_440_1279 = not_525_1109 ^ not_403_1234;
assign not_450_1280 = ~xor_450_1279;
assign xor_450_1279 = gate3_357_1182 ^ xor_435_1233;
assign gate3_317_1366 = xor_440_1279 & gate3_306_1330;
assign xor_314_1394 = not_306_1367 ^ not_422_1280;
assign gate3_243_1453 = xor_314_1394 | not_244_1452;
assign not_244_1452 = ~gate3_238_1430;
assign xor_217_1478 = xor_305_1394 ^ xor_237_1453;
assign gate3_241_1430 = gate3_323_1366 & gate3_319_1394;
assign gate3_319_1394 = gate3_363_1182 | xor_326_1366;
assign gate3_323_1366 = not_456_1280 | not_324_1365;
assign not_324_1365 = ~gate3_309_1330;
assign gate3_150_1576 = gate3_191_1528 | gate3_187_1555;
assign gate3_187_1555 = gate3_247_1430 & not_194_1529;
assign not_194_1529 = ~xor_194_1528;
assign xor_194_1528 = xor_231_1478 ^ gate3_167_1503;
assign gate3_167_1503 = gate3_252_1453 & gate3_223_1478;
assign gate3_223_1478 = xor_346_1394 | xor_255_1453;
assign xor_255_1453 = gate3_244_1430 ^ not_337_1395;
assign not_337_1395 = ~xor_337_1394;
assign xor_337_1394 = not_450_1280 ^ xor_320_1366;
assign gate3_244_1430 = gate3_329_1366 | gate3_331_1394;
assign gate3_331_1394 = not_332_1393 & not_475_1280;
assign not_475_1280 = ~xor_475_1279;
assign xor_475_1279 = gate3_369_1182 ^ not_451_1234;
assign not_451_1234 = ~xor_451_1233;
assign xor_451_1233 = xor_597_1108 ^ gate3_374_1182;
assign gate3_374_1182 = gate3_586_1108 & gate3_584_1054;
assign gate3_584_1054 = not_876_858 | not_585_1053;
assign not_585_1053 = ~gate3_477_983;
assign gate3_477_983 = gate3_1006_774 | gate3_861_857;
assign gate3_861_857 = gate3_1046_728 & xor_1009_774;
assign xor_1009_774 = gate3_1004_728 ^ gate3_1049_728;
assign gate3_1049_728 = lever[24] & lever[10];
assign gate3_1004_728 = lever[23] & lever[11];
assign gate3_1046_728 = lever[25] & lever[9];
assign gate3_1006_774 = gate3_1004_728 & gate3_1049_728;
assign not_876_858 = ~xor_876_857;
assign xor_876_857 = gate3_1013_728 ^ xor_961_774;
assign gate3_586_1108 = xor_589_1054 | not_587_1107;
assign not_587_1107 = ~gate3_474_983;
assign gate3_474_983 = gate3_1015_774 | gate3_873_857;
assign gate3_873_857 = xor_1018_774 & gate3_1061_728;
assign gate3_1061_728 = lever[6] & lever[28];
assign xor_1018_774 = gate3_1010_728 ^ gate3_1055_728;
assign gate3_1055_728 = lever[7] & lever[27];
assign gate3_1010_728 = lever[8] & lever[26];
assign gate3_1015_774 = gate3_1010_728 & gate3_1055_728;
assign xor_589_1054 = not_876_858 ^ gate3_477_983;
assign xor_597_1108 = not_846_858 ^ xor_569_1054;
assign gate3_369_1182 = gate3_592_1054 & gate3_594_1108;
assign gate3_594_1108 = xor_595_1054 | not_888_858;
assign not_888_858 = ~xor_888_857;
assign xor_888_857 = gate3_1031_728 ^ xor_991_774;
assign xor_595_1054 = gate3_482_983 ^ not_882_858;
assign not_882_858 = ~xor_882_857;
assign xor_882_857 = gate3_1022_728 ^ xor_970_774;
assign gate3_482_983 = gate3_1024_774 | gate3_879_857;
assign gate3_879_857 = xor_1027_774 & gate3_1070_728;
assign gate3_1070_728 = lever[3] & lever[31];
assign xor_1027_774 = gate3_1019_728 ^ gate3_1064_728;
assign gate3_1064_728 = lever[30] & lever[4];
assign gate3_1019_728 = lever[29] & lever[5];
assign gate3_1024_774 = gate3_1019_728 & gate3_1064_728;
assign gate3_592_1054 = not_882_858 | not_593_1053;
assign not_593_1053 = ~gate3_482_983;
assign not_332_1393 = ~not_332_1367;
assign not_332_1367 = ~xor_332_1366;
assign xor_332_1366 = not_468_1280 ^ gate3_312_1330;
assign gate3_312_1330 = gate3_438_1233 | gate3_462_1279;
assign gate3_462_1279 = not_441_1234 & not_589_1109;
assign not_589_1109 = ~xor_589_1108;
assign xor_589_1108 = gate3_474_983 ^ xor_589_1054;
assign not_441_1234 = ~xor_441_1233;
assign xor_441_1233 = xor_580_1108 ^ gate3_366_1182;
assign gate3_366_1182 = gate3_578_1054 & gate3_570_1108;
assign gate3_570_1108 = not_867_858 | xor_581_1054;
assign xor_581_1054 = not_858_858 ^ gate3_471_983;
assign gate3_471_983 = gate3_1000_774 | gate3_852_857;
assign gate3_852_857 = gate3_1043_728 & xor_1003_774;
assign xor_1003_774 = gate3_992_728 ^ gate3_1037_728;
assign gate3_1037_728 = lever[12] & lever[21];
assign gate3_992_728 = lever[13] & lever[20];
assign gate3_1043_728 = lever[22] & lever[11];
assign gate3_1000_774 = gate3_992_728 & gate3_1037_728;
assign not_858_858 = ~xor_858_857;
assign xor_858_857 = gate3_995_728 ^ xor_946_774;
assign not_867_858 = ~xor_867_857;
assign xor_867_857 = gate3_1046_728 ^ xor_1009_774;
assign gate3_578_1054 = not_858_858 | not_579_1053;
assign not_579_1053 = ~gate3_471_983;
assign xor_580_1108 = not_822_858 ^ xor_551_1054;
assign gate3_438_1233 = xor_580_1108 & not_439_1232;
assign not_439_1232 = ~gate3_366_1182;
assign not_468_1280 = ~xor_468_1279;
assign xor_468_1279 = xor_558_1108 ^ not_429_1234;
assign gate3_329_1366 = not_468_1280 & gate3_312_1330;
assign xor_346_1394 = xor_338_1366 ^ gate3_600_1108;
assign gate3_600_1108 = gate3_598_1054 & xor_601_1054;
assign xor_601_1054 = xor_976_774 ^ gate3_467_983;
assign gate3_598_1054 = gate3_980_728 & gate3_485_983;
assign gate3_485_983 = gate3_1036_774 | gate3_894_857;
assign gate3_894_857 = gate3_1079_728 & xor_1039_774;
assign xor_1039_774 = gate3_1073_728 ^ gate3_1028_728;
assign gate3_1028_728 = lever[2] & lever[32];
assign gate3_1073_728 = lever[1] & lever[33];
assign gate3_1079_728 = lever[34] & lever[0];
assign gate3_1036_774 = gate3_1028_728 & gate3_1073_728;
assign xor_338_1366 = xor_377_1182 ^ gate3_317_1330;
assign gate3_317_1330 = gate3_448_1233 | gate3_471_1279;
assign gate3_471_1279 = not_451_1234 & not_472_1278;
assign not_472_1278 = ~gate3_369_1182;
assign gate3_448_1233 = xor_597_1108 & not_449_1232;
assign not_449_1232 = ~gate3_374_1182;
assign xor_377_1182 = xor_575_1054 ^ gate3_603_1108;
assign gate3_603_1108 = gate3_934_774 | gate3_572_1054;
assign gate3_252_1453 = not_337_1395 | not_253_1452;
assign not_253_1452 = ~gate3_244_1430;
assign xor_231_1478 = not_325_1395 ^ xor_249_1453;
assign gate3_247_1430 = gate3_335_1366 | gate3_343_1394;
assign gate3_343_1394 = gate3_600_1108 & not_344_1393;
assign not_344_1393 = ~xor_338_1366;
assign gate3_335_1366 = gate3_317_1330 & not_336_1365;
assign not_336_1365 = ~xor_377_1182;
assign gate3_191_1528 = xor_231_1478 & not_192_1527;
assign not_192_1527 = ~gate3_167_1503;
assign gate3_180_1628 = gate3_1082_728 & not_181_1627;
assign not_181_1627 = ~not_165_1603;
assign not_165_1603 = ~xor_165_1602;
assign xor_165_1602 = gate3_150_1576 ^ not_193_1556;
assign gate3_1082_728 = lever[0] & lever[39];
assign not_183_1629 = ~xor_183_1628;
assign xor_183_1628 = gate3_1034_728 ^ xor_159_1602;
assign xor_159_1602 = not_181_1556 ^ gate3_147_1576;
assign gate3_147_1576 = gate3_185_1528 | not_148_1575;
assign not_148_1575 = ~gate3_175_1555;
assign gate3_175_1555 = not_176_1554 | gate3_241_1430;
assign not_176_1554 = ~not_188_1529;
assign gate3_185_1528 = xor_217_1478 & not_186_1527;
assign not_186_1527 = ~gate3_164_1503;
assign not_181_1556 = ~xor_181_1555;
assign xor_181_1555 = gate3_235_1430 ^ xor_182_1528;
assign gate3_1034_728 = lever[1] & lever[39];
assign xor_43_1679 = gate3_141_1654 ^ not_177_1629;
assign not_177_1629 = ~xor_177_1628;
assign xor_177_1628 = gate3_986_728 ^ not_153_1603;
assign gate3_141_1654 = gate3_167_1628 | gate3_156_1602;
assign gate3_156_1602 = gate3_147_1576 & not_181_1556;
assign gate3_167_1628 = xor_159_1602 & gate3_1034_728;
assign gate3_49_1679 = not_177_1629 | not_50_1678;
assign not_50_1678 = ~gate3_141_1654;
assign gate3_1_1800 = gate3_1_1793 | xor_43_1679;
assign gate3_1_1793 = gate3_1_1785 | xor_11_1679;
assign xor_11_1679 = gate3_144_1654 ^ not_183_1629;
assign gate3_1_1785 = gate3_1_1778 & gate3_39_1654;
assign gate3_39_1654 = gate3_169_1602 | xor_186_1628;
assign xor_186_1628 = gate3_1082_728 ^ not_165_1603;
assign gate3_169_1602 = not_205_1556 | not_170_1601;
assign not_170_1601 = ~gate3_153_1576;
assign gate3_153_1576 = gate3_197_1528 | not_154_1575;
assign not_154_1575 = ~gate3_199_1555;
assign gate3_199_1555 = gate3_349_1366 | not_200_1554;
assign not_200_1554 = ~not_200_1529;
assign not_200_1529 = ~xor_200_1528;
assign xor_200_1528 = gate3_170_1503 ^ xor_245_1478;
assign xor_245_1478 = xor_346_1394 ^ xor_255_1453;
assign gate3_170_1503 = gate3_261_1453 & gate3_237_1478;
assign gate3_237_1478 = xor_352_1366 | xor_264_1453;
assign xor_264_1453 = gate3_253_1430 ^ xor_360_1394;
assign xor_360_1394 = not_475_1280 ^ not_332_1367;
assign gate3_253_1430 = gate3_341_1366 | gate3_357_1394;
assign gate3_357_1394 = not_505_1280 & not_358_1393;
assign not_358_1393 = ~not_344_1367;
assign not_344_1367 = ~xor_344_1366;
assign xor_344_1366 = gate3_320_1330 ^ xor_487_1279;
assign xor_487_1279 = not_589_1109 ^ not_441_1234;
assign gate3_320_1330 = gate3_454_1233 | gate3_481_1279;
assign gate3_481_1279 = not_621_1109 & not_457_1234;
assign not_457_1234 = ~xor_457_1233;
assign xor_457_1233 = xor_610_1108 ^ gate3_380_1182;
assign gate3_380_1182 = gate3_605_1054 & gate3_607_1108;
assign gate3_607_1108 = xor_608_1054 | not_912_858;
assign not_912_858 = ~xor_912_857;
assign xor_912_857 = gate3_1094_728 ^ xor_1057_774;
assign xor_1057_774 = gate3_1097_728 ^ gate3_1052_728;
assign gate3_1052_728 = lever[23] & lever[10];
assign gate3_1097_728 = lever[9] & lever[24];
assign gate3_1094_728 = lever[8] & lever[25];
assign xor_608_1054 = gate3_491_983 ^ not_903_858;
assign not_903_858 = ~xor_903_857;
assign xor_903_857 = gate3_1043_728 ^ xor_1003_774;
assign gate3_491_983 = gate3_1048_774 | gate3_900_857;
assign gate3_900_857 = gate3_1091_728 & xor_1051_774;
assign xor_1051_774 = gate3_1040_728 ^ gate3_1085_728;
assign gate3_1085_728 = lever[11] & lever[21];
assign gate3_1040_728 = lever[12] & lever[20];
assign gate3_1091_728 = lever[22] & lever[10];
assign gate3_1048_774 = gate3_1040_728 & gate3_1085_728;
assign gate3_605_1054 = not_903_858 | not_606_1053;
assign not_606_1053 = ~gate3_491_983;
assign xor_610_1108 = not_867_858 ^ xor_581_1054;
assign not_621_1109 = ~xor_621_1108;
assign xor_621_1108 = gate3_494_983 ^ xor_621_1054;
assign xor_621_1054 = not_931_858 ^ gate3_497_983;
assign gate3_497_983 = gate3_1054_774 | gate3_909_857;
assign gate3_909_857 = gate3_1094_728 & xor_1057_774;
assign gate3_1054_774 = gate3_1052_728 & gate3_1097_728;
assign not_931_858 = ~xor_931_857;
assign xor_931_857 = xor_1018_774 ^ gate3_1061_728;
assign gate3_494_983 = gate3_1063_774 | gate3_915_857;
assign gate3_915_857 = gate3_1109_728 & xor_1066_774;
assign xor_1066_774 = gate3_1058_728 ^ gate3_1103_728;
assign gate3_1103_728 = lever[6] & lever[27];
assign gate3_1058_728 = lever[26] & lever[7];
assign gate3_1109_728 = lever[5] & lever[28];
assign gate3_1063_774 = gate3_1055_728 & gate3_1106_728;
assign gate3_1106_728 = lever[26] & lever[6];
assign gate3_454_1233 = xor_610_1108 & not_455_1232;
assign not_455_1232 = ~gate3_380_1182;
assign not_505_1280 = ~xor_505_1279;
assign xor_505_1279 = gate3_384_1182 ^ not_463_1234;
assign not_463_1234 = ~xor_463_1233;
assign xor_463_1233 = xor_632_1108 ^ gate3_389_1182;
assign gate3_389_1182 = gate3_614_1054 & gate3_616_1108;
assign gate3_616_1108 = not_617_1107 | xor_621_1054;
assign not_617_1107 = ~gate3_494_983;
assign gate3_614_1054 = not_931_858 | not_615_1053;
assign not_615_1053 = ~gate3_497_983;
assign xor_632_1108 = not_888_858 ^ xor_595_1054;
assign gate3_384_1182 = gate3_624_1054 & gate3_626_1108;
assign gate3_626_1108 = not_945_858 | xor_627_1054;
assign xor_627_1054 = gate3_503_983 ^ not_939_858;
assign not_939_858 = ~xor_939_857;
assign xor_939_857 = gate3_1070_728 ^ xor_1027_774;
assign gate3_503_983 = gate3_1072_774 | gate3_936_857;
assign gate3_936_857 = xor_1075_774 & gate3_1118_728;
assign gate3_1118_728 = lever[2] & lever[31];
assign xor_1075_774 = gate3_1067_728 ^ gate3_1112_728;
assign gate3_1112_728 = lever[3] & lever[30];
assign gate3_1067_728 = lever[29] & lever[4];
assign gate3_1072_774 = gate3_1067_728 & gate3_1112_728;
assign not_945_858 = ~xor_945_857;
assign xor_945_857 = gate3_1079_728 ^ xor_1039_774;
assign gate3_624_1054 = not_939_858 | not_625_1053;
assign not_625_1053 = ~gate3_503_983;
assign gate3_341_1366 = gate3_320_1330 & xor_487_1279;
assign xor_352_1366 = gate3_326_1330 ^ not_638_1109;
assign not_638_1109 = ~xor_638_1108;
assign xor_638_1108 = gate3_598_1054 ^ xor_601_1054;
assign gate3_326_1330 = gate3_460_1233 | gate3_496_1279;
assign gate3_496_1279 = not_463_1234 & not_497_1278;
assign not_497_1278 = ~gate3_384_1182;
assign gate3_460_1233 = not_461_1232 & xor_632_1108;
assign not_461_1232 = ~gate3_389_1182;
assign gate3_261_1453 = xor_360_1394 | not_262_1452;
assign not_262_1452 = ~gate3_253_1430;
assign gate3_349_1366 = not_638_1109 | not_350_1365;
assign not_350_1365 = ~gate3_326_1330;
assign gate3_197_1528 = xor_245_1478 & not_198_1527;
assign not_198_1527 = ~gate3_170_1503;
assign not_205_1556 = ~xor_205_1555;
assign xor_205_1555 = gate3_247_1430 ^ not_194_1529;
assign gate3_1_1778 = gate3_1_1770 | not_14_1655;
assign not_14_1655 = ~xor_14_1654;
assign xor_14_1654 = gate3_169_1602 ^ xor_186_1628;
assign gate3_1_1770 = gate3_1_1764 & gate3_9_1654;
assign gate3_9_1654 = not_172_1628 | xor_175_1602;
assign xor_175_1602 = gate3_153_1576 ^ not_205_1556;
assign not_172_1628 = ~gate3_172_1602;
assign gate3_172_1602 = not_211_1556 & gate3_158_1576;
assign gate3_158_1576 = gate3_203_1528 | gate3_208_1555;
assign gate3_208_1555 = not_206_1529 & gate3_365_1366;
assign gate3_365_1366 = xor_648_1054 & gate3_332_1330;
assign gate3_332_1330 = gate3_473_1233 | gate3_520_1279;
assign gate3_520_1279 = not_476_1234 & not_521_1278;
assign not_521_1278 = ~gate3_398_1182;
assign gate3_398_1182 = gate3_642_1054 & gate3_672_1108;
assign gate3_672_1108 = not_1123_775 | xor_645_1054;
assign xor_645_1054 = not_990_858 ^ gate3_529_983;
assign gate3_529_983 = gate3_1111_774 | gate3_978_857;
assign gate3_978_857 = gate3_1154_728 & xor_1114_774;
assign xor_1114_774 = gate3_1115_728 ^ gate3_1148_728;
assign gate3_1148_728 = lever[2] & lever[30];
assign gate3_1115_728 = lever[29] & lever[3];
assign gate3_1154_728 = lever[1] & lever[31];
assign gate3_1111_774 = gate3_1115_728 & gate3_1148_728;
assign not_990_858 = ~xor_990_857;
assign xor_990_857 = gate3_1118_728 ^ xor_1075_774;
assign not_1123_775 = ~xor_1123_774;
assign xor_1123_774 = gate3_1076_728 ^ gate3_1157_728;
assign gate3_1157_728 = lever[0] & lever[33];
assign gate3_1076_728 = lever[1] & lever[32];
assign gate3_642_1054 = not_643_1053 | not_990_858;
assign not_643_1053 = ~gate3_529_983;
assign not_476_1234 = ~xor_476_1233;
assign xor_476_1233 = xor_681_1108 ^ gate3_403_1182;
assign gate3_403_1182 = gate3_636_1054 & gate3_663_1108;
assign gate3_663_1108 = xor_639_1054 | not_664_1107;
assign not_664_1107 = ~gate3_512_983;
assign gate3_512_983 = gate3_1102_774 | gate3_969_857;
assign gate3_969_857 = gate3_1145_728 & xor_1105_774;
assign xor_1105_774 = gate3_1139_728 ^ gate3_1106_728;
assign gate3_1139_728 = lever[27] & lever[5];
assign gate3_1145_728 = lever[4] & lever[28];
assign gate3_1102_774 = gate3_1106_728 & gate3_1139_728;
assign xor_639_1054 = not_972_858 ^ gate3_518_983;
assign gate3_518_983 = gate3_1096_774 | gate3_960_857;
assign gate3_960_857 = xor_1099_774 & gate3_1130_728;
assign gate3_1130_728 = lever[25] & lever[7];
assign xor_1099_774 = gate3_1133_728 ^ gate3_1100_728;
assign gate3_1100_728 = lever[23] & lever[9];
assign gate3_1133_728 = lever[24] & lever[8];
assign gate3_1096_774 = gate3_1100_728 & gate3_1133_728;
assign not_972_858 = ~xor_972_857;
assign xor_972_857 = gate3_1109_728 ^ xor_1066_774;
assign gate3_636_1054 = not_972_858 | not_637_1053;
assign not_637_1053 = ~gate3_518_983;
assign xor_681_1108 = not_945_858 ^ xor_627_1054;
assign gate3_473_1233 = xor_681_1108 & not_474_1232;
assign not_474_1232 = ~gate3_403_1182;
assign xor_648_1054 = gate3_980_728 ^ gate3_485_983;
assign not_206_1529 = ~xor_206_1528;
assign xor_206_1528 = xor_254_1478 ^ gate3_173_1503;
assign gate3_173_1503 = gate3_249_1478 & gate3_270_1453;
assign gate3_270_1453 = xor_373_1394 | not_271_1452;
assign not_271_1452 = ~gate3_256_1430;
assign gate3_256_1430 = gate3_355_1366 | gate3_363_1394;
assign gate3_363_1394 = not_364_1393 & not_523_1280;
assign not_523_1280 = ~xor_523_1279;
assign xor_523_1279 = gate3_398_1182 ^ not_476_1234;
assign not_364_1393 = ~not_359_1367;
assign not_359_1367 = ~xor_359_1366;
assign xor_359_1366 = gate3_329_1330 ^ xor_517_1279;
assign xor_517_1279 = not_621_1109 ^ not_457_1234;
assign gate3_329_1330 = gate3_466_1233 | gate3_514_1279;
assign gate3_514_1279 = not_666_1109 & not_469_1234;
assign not_469_1234 = ~xor_469_1233;
assign xor_469_1233 = gate3_393_1182 ^ xor_658_1108;
assign xor_658_1108 = not_912_858 ^ xor_608_1054;
assign gate3_393_1182 = gate3_630_1054 & gate3_644_1108;
assign gate3_644_1108 = not_963_858 | xor_633_1054;
assign xor_633_1054 = gate3_509_983 ^ not_954_858;
assign not_954_858 = ~xor_954_857;
assign xor_954_857 = gate3_1091_728 ^ xor_1051_774;
assign gate3_509_983 = gate3_1084_774 | gate3_951_857;
assign gate3_951_857 = gate3_1127_728 & xor_1087_774;
assign xor_1087_774 = gate3_1088_728 ^ gate3_1121_728;
assign gate3_1121_728 = lever[10] & lever[21];
assign gate3_1088_728 = lever[20] & lever[11];
assign gate3_1127_728 = lever[22] & lever[9];
assign gate3_1084_774 = gate3_1088_728 & gate3_1121_728;
assign not_963_858 = ~xor_963_857;
assign xor_963_857 = gate3_1130_728 ^ xor_1099_774;
assign gate3_630_1054 = not_954_858 | not_631_1053;
assign not_631_1053 = ~gate3_509_983;
assign not_666_1109 = ~xor_666_1108;
assign xor_666_1108 = gate3_512_983 ^ xor_639_1054;
assign gate3_466_1233 = xor_658_1108 & not_467_1232;
assign not_467_1232 = ~gate3_393_1182;
assign gate3_355_1366 = gate3_329_1330 & xor_517_1279;
assign xor_373_1394 = not_505_1280 ^ not_344_1367;
assign gate3_249_1478 = not_368_1367 | xor_273_1453;
assign xor_273_1453 = gate3_256_1430 ^ xor_373_1394;
assign not_368_1367 = ~xor_368_1366;
assign xor_368_1366 = xor_648_1054 ^ gate3_332_1330;
assign xor_254_1478 = xor_352_1366 ^ xor_264_1453;
assign gate3_203_1528 = xor_254_1478 & not_204_1527;
assign not_204_1527 = ~gate3_173_1503;
assign not_211_1556 = ~xor_211_1555;
assign xor_211_1555 = gate3_349_1366 ^ not_200_1529;
assign gate3_1_1764 = gate3_1_1756 | xor_41_1628;
assign xor_41_1628 = gate3_172_1602 ^ xor_175_1602;
assign gate3_1_1756 = gate3_1_1749 | gate3_37_1628;
assign gate3_37_1628 = not_181_1603 & gate3_178_1602;
assign gate3_178_1602 = gate3_164_1576 | not_219_1556;
assign not_219_1556 = ~xor_219_1555;
assign xor_219_1555 = gate3_365_1366 ^ not_206_1529;
assign gate3_164_1576 = gate3_214_1528 & not_165_1575;
assign not_165_1575 = ~gate3_216_1555;
assign gate3_216_1555 = gate3_377_1366 & xor_217_1528;
assign xor_217_1528 = gate3_176_1503 ^ not_263_1479;
assign not_263_1479 = ~xor_263_1478;
assign xor_263_1478 = not_368_1367 ^ xor_273_1453;
assign gate3_176_1503 = gate3_276_1453 & gate3_257_1478;
assign gate3_257_1478 = xor_380_1366 | xor_279_1453;
assign xor_279_1453 = gate3_261_1430 ^ xor_394_1394;
assign xor_394_1394 = not_523_1280 ^ not_359_1367;
assign gate3_261_1430 = gate3_371_1366 | gate3_391_1394;
assign gate3_391_1394 = xor_535_1279 & xor_374_1366;
assign xor_374_1366 = xor_529_1279 ^ gate3_335_1330;
assign gate3_335_1330 = gate3_479_1233 | not_336_1329;
assign not_336_1329 = ~gate3_526_1279;
assign gate3_526_1279 = xor_709_1108 | not_527_1278;
assign not_527_1278 = ~not_482_1234;
assign not_482_1234 = ~xor_482_1233;
assign xor_482_1233 = xor_702_1108 ^ gate3_406_1182;
assign gate3_406_1182 = gate3_684_1108 & gate3_651_1054;
assign gate3_651_1054 = not_996_858 | not_652_1053;
assign not_652_1053 = ~gate3_533_983;
assign gate3_533_983 = gate3_1132_774 | gate3_993_857;
assign gate3_993_857 = gate3_1169_728 & xor_1135_774;
assign xor_1135_774 = gate3_1124_728 ^ gate3_1163_728;
assign gate3_1163_728 = lever[21] & lever[9];
assign gate3_1124_728 = lever[10] & lever[20];
assign gate3_1169_728 = lever[22] & lever[8];
assign gate3_1132_774 = gate3_1124_728 & gate3_1163_728;
assign not_996_858 = ~xor_996_857;
assign xor_996_857 = gate3_1127_728 ^ xor_1087_774;
assign gate3_684_1108 = not_1008_858 | xor_658_1054;
assign xor_658_1054 = gate3_533_983 ^ not_996_858;
assign not_1008_858 = ~xor_1008_857;
assign xor_1008_857 = gate3_1172_728 ^ xor_1141_774;
assign xor_1141_774 = gate3_1136_728 ^ gate3_1175_728;
assign gate3_1175_728 = lever[24] & lever[7];
assign gate3_1136_728 = lever[23] & lever[8];
assign gate3_1172_728 = lever[25] & lever[6];
assign xor_702_1108 = not_963_858 ^ xor_633_1054;
assign xor_709_1108 = gate3_536_983 ^ xor_665_1054;
assign xor_665_1054 = not_1017_858 ^ gate3_539_983;
assign gate3_539_983 = gate3_1138_774 | gate3_1002_857;
assign gate3_1002_857 = gate3_1172_728 & xor_1141_774;
assign gate3_1138_774 = gate3_1136_728 & gate3_1175_728;
assign not_1017_858 = ~xor_1017_857;
assign xor_1017_857 = gate3_1145_728 ^ xor_1105_774;
assign gate3_536_983 = gate3_1147_774 | gate3_1011_857;
assign gate3_1011_857 = gate3_1187_728 & xor_1150_774;
assign xor_1150_774 = gate3_1142_728 ^ gate3_1181_728;
assign gate3_1181_728 = lever[4] & lever[27];
assign gate3_1142_728 = lever[26] & lever[5];
assign gate3_1187_728 = lever[3] & lever[28];
assign gate3_1147_774 = gate3_1142_728 & gate3_1181_728;
assign gate3_479_1233 = xor_702_1108 & not_480_1232;
assign not_480_1232 = ~gate3_406_1182;
assign xor_529_1279 = not_666_1109 ^ not_469_1234;
assign xor_535_1279 = gate3_409_1182 ^ not_488_1234;
assign not_488_1234 = ~xor_488_1233;
assign xor_488_1233 = gate3_414_1182 ^ not_718_1109;
assign not_718_1109 = ~xor_718_1108;
assign xor_718_1108 = not_1123_775 ^ xor_645_1054;
assign gate3_414_1182 = gate3_661_1054 & gate3_705_1108;
assign gate3_705_1108 = xor_665_1054 | not_706_1107;
assign not_706_1107 = ~gate3_536_983;
assign gate3_661_1054 = not_1017_858 | not_662_1053;
assign not_662_1053 = ~gate3_539_983;
assign gate3_409_1182 = gate3_670_1054 & not_410_1181;
assign not_410_1181 = ~gate3_712_1108;
assign gate3_712_1108 = gate3_1160_728 & not_713_1107;
assign not_713_1107 = ~xor_673_1054;
assign xor_673_1054 = not_1026_858 ^ gate3_545_983;
assign gate3_545_983 = gate3_1156_774 | gate3_1020_857;
assign gate3_1020_857 = gate3_1196_728 & xor_1162_774;
assign xor_1162_774 = gate3_1190_728 ^ gate3_1151_728;
assign gate3_1151_728 = lever[29] & lever[2];
assign gate3_1190_728 = lever[30] & lever[1];
assign gate3_1196_728 = lever[0] & lever[31];
assign gate3_1156_774 = gate3_1151_728 & gate3_1190_728;
assign not_1026_858 = ~xor_1026_857;
assign xor_1026_857 = gate3_1154_728 ^ xor_1114_774;
assign gate3_1160_728 = lever[0] & lever[32];
assign gate3_670_1054 = not_1026_858 | not_671_1053;
assign not_671_1053 = ~gate3_545_983;
assign gate3_371_1366 = xor_529_1279 & gate3_335_1330;
assign xor_380_1366 = gate3_1120_774 ^ gate3_340_1330;
assign gate3_340_1330 = gate3_485_1233 & gate3_532_1279;
assign gate3_532_1279 = gate3_409_1182 | not_488_1234;
assign gate3_485_1233 = gate3_414_1182 | not_718_1109;
assign gate3_1120_774 = gate3_1073_728 & gate3_1160_728;
assign gate3_276_1453 = xor_394_1394 | not_277_1452;
assign not_277_1452 = ~gate3_261_1430;
assign gate3_377_1366 = gate3_1120_774 & not_378_1365;
assign not_378_1365 = ~gate3_340_1330;
assign gate3_214_1528 = gate3_176_1503 | not_263_1479;
assign not_181_1603 = ~xor_181_1602;
assign xor_181_1602 = gate3_158_1576 ^ not_211_1556;
assign gate3_1_1749 = gate3_1_1743 & gate3_34_1628;
assign gate3_34_1628 = gate3_178_1602 | not_181_1603;
assign gate3_1_1743 = gate3_1_1736 | gate3_28_1628;
assign gate3_28_1628 = gate3_167_1576 & not_29_1627;
assign not_29_1627 = ~xor_184_1602;
assign xor_184_1602 = not_219_1556 ^ gate3_164_1576;
assign gate3_167_1576 = gate3_51_1528 | not_37_1556;
assign not_37_1556 = ~xor_37_1555;
assign xor_37_1555 = gate3_377_1366 ^ xor_217_1528;
assign gate3_51_1528 = not_47_1479 | gate3_36_1503;
assign gate3_36_1503 = gate3_285_1453 & gate3_266_1478;
assign gate3_266_1478 = gate3_51_1330 | xor_45_1453;
assign xor_45_1453 = gate3_264_1430 ^ not_400_1395;
assign not_400_1395 = ~xor_400_1394;
assign xor_400_1394 = xor_535_1279 ^ xor_374_1366;
assign gate3_264_1430 = gate3_383_1366 | gate3_397_1394;
assign gate3_397_1394 = xor_25_1279 & xor_23_1366;
assign xor_23_1366 = gate3_343_1330 ^ not_541_1280;
assign not_541_1280 = ~xor_541_1279;
assign xor_541_1279 = xor_709_1108 ^ not_482_1234;
assign gate3_343_1330 = gate3_491_1233 | not_344_1329;
assign not_344_1329 = ~gate3_538_1279;
assign gate3_538_1279 = not_539_1278 | xor_24_1108;
assign xor_24_1108 = gate3_554_983 ^ xor_682_1054;
assign xor_682_1054 = not_1044_858 ^ gate3_557_983;
assign gate3_557_983 = gate3_1038_857 | gate3_1177_774;
assign gate3_1177_774 = gate3_1178_728 & gate3_1211_728;
assign gate3_1211_728 = lever[6] & lever[24];
assign gate3_1178_728 = lever[23] & lever[7];
assign gate3_1038_857 = gate3_1208_728 & xor_1180_774;
assign xor_1180_774 = gate3_1211_728 ^ gate3_1178_728;
assign gate3_1208_728 = lever[5] & lever[25];
assign not_1044_858 = ~xor_1044_857;
assign xor_1044_857 = gate3_1187_728 ^ xor_1150_774;
assign gate3_554_983 = gate3_1041_857 | gate3_1183_774;
assign gate3_1183_774 = gate3_1184_728 & gate3_1217_728;
assign gate3_1217_728 = lever[27] & lever[3];
assign gate3_1184_728 = lever[4] & lever[26];
assign gate3_1041_857 = xor_1192_774 & gate3_1223_728;
assign gate3_1223_728 = lever[2] & lever[28];
assign xor_1192_774 = gate3_1184_728 ^ gate3_1217_728;
assign not_539_1278 = ~not_22_1234;
assign not_22_1234 = ~xor_22_1233;
assign xor_22_1233 = gate3_417_1182 ^ xor_727_1108;
assign xor_727_1108 = not_1008_858 ^ xor_658_1054;
assign gate3_417_1182 = gate3_676_1054 & gate3_724_1108;
assign gate3_724_1108 = not_3_858 | xor_13_1054;
assign xor_13_1054 = gate3_548_983 ^ not_1032_858;
assign not_1032_858 = ~xor_1032_857;
assign xor_1032_857 = xor_1135_774 ^ gate3_1169_728;
assign gate3_548_983 = gate3_1029_857 | gate3_1165_774;
assign gate3_1165_774 = gate3_1166_728 & gate3_1199_728;
assign gate3_1199_728 = lever[21] & lever[8];
assign gate3_1166_728 = lever[20] & lever[9];
assign gate3_1029_857 = gate3_1205_728 & xor_1174_774;
assign xor_1174_774 = gate3_1166_728 ^ gate3_1199_728;
assign gate3_1205_728 = lever[22] & lever[7];
assign not_3_858 = ~xor_3_857;
assign xor_3_857 = gate3_1208_728 ^ xor_1180_774;
assign gate3_676_1054 = not_1032_858 | not_677_1053;
assign not_677_1053 = ~gate3_548_983;
assign gate3_491_1233 = xor_727_1108 & not_492_1232;
assign not_492_1232 = ~gate3_417_1182;
assign xor_25_1279 = gate3_560_983 ^ not_497_1234;
assign not_497_1234 = ~xor_497_1233;
assign xor_497_1233 = xor_733_1108 ^ gate3_424_1182;
assign gate3_424_1182 = gate3_679_1054 & gate3_730_1108;
assign gate3_730_1108 = not_731_1107 | xor_682_1054;
assign not_731_1107 = ~gate3_554_983;
assign gate3_679_1054 = not_1044_858 | not_680_1053;
assign not_680_1053 = ~gate3_557_983;
assign xor_733_1108 = gate3_1160_728 ^ xor_673_1054;
assign gate3_560_983 = gate3_6_857 | not_9_858;
assign not_9_858 = ~xor_9_857;
assign xor_9_857 = gate3_1196_728 ^ xor_1162_774;
assign gate3_6_857 = not_1190_774 | not_7_856;
assign not_7_856 = ~gate3_1229_728;
assign gate3_1229_728 = lever[0] & lever[29];
assign not_1190_774 = ~gate3_1190_728;
assign gate3_383_1366 = gate3_343_1330 & not_541_1280;
assign gate3_51_1330 = gate3_494_1233 & gate3_544_1279;
assign gate3_544_1279 = gate3_560_983 | not_497_1234;
assign gate3_494_1233 = xor_733_1108 | gate3_424_1182;
assign gate3_285_1453 = not_400_1395 | not_286_1452;
assign not_286_1452 = ~gate3_264_1430;
assign not_47_1479 = ~xor_47_1478;
assign xor_47_1478 = xor_380_1366 ^ xor_279_1453;
assign gate3_1_1736 = not_2_1735 & gate3_25_1628;
assign gate3_25_1628 = not_26_1627 | gate3_167_1576;
assign not_26_1627 = ~xor_184_1602;
assign not_2_1735 = ~gate3_1_1728;
assign gate3_1_1728 = not_2_1727 | gate3_22_1628;
assign gate3_22_1628 = gate3_20_1602 | gate3_32_1602;
assign gate3_32_1602 = xor_24_1576 & gate3_30_1576;
assign gate3_30_1576 = gate3_17_1555 & not_31_1575;
assign not_31_1575 = ~not_40_1556;
assign not_40_1556 = ~xor_40_1555;
assign xor_40_1555 = xor_45_1528 ^ gate3_38_1528;
assign gate3_38_1528 = not_39_1527 & xor_44_1478;
assign xor_44_1478 = xor_45_1453 ^ gate3_51_1330;
assign not_39_1527 = ~gate3_33_1503;
assign gate3_33_1503 = gate3_20_1453 & gate3_22_1478;
assign gate3_22_1478 = xor_23_1453 | gate3_15_1233;
assign gate3_15_1233 = gate3_7_1182 | not_5_984;
assign not_5_984 = ~xor_5_983;
assign xor_5_983 = gate3_6_857 ^ not_9_858;
assign gate3_7_1182 = gate3_16_1054 & gate3_21_1108;
assign gate3_21_1108 = xor_7_1054 | not_22_1107;
assign not_22_1107 = ~gate3_1_983;
assign gate3_1_983 = gate3_1113_857 | gate3_1273_774;
assign gate3_1273_774 = gate3_1220_728 & gate3_1295_728;
assign gate3_1295_728 = lever[27] & lever[2];
assign gate3_1220_728 = lever[26] & lever[3];
assign gate3_1113_857 = gate3_1310_728 & xor_1276_774;
assign xor_1276_774 = gate3_1220_728 ^ gate3_1295_728;
assign gate3_1310_728 = lever[1] & lever[28];
assign xor_7_1054 = gate3_599_983 ^ not_1140_858;
assign not_1140_858 = ~xor_1140_857;
assign xor_1140_857 = gate3_1223_728 ^ xor_1192_774;
assign gate3_599_983 = gate3_1279_774 | gate3_1125_857;
assign gate3_1125_857 = xor_1282_774 & gate3_1313_728;
assign gate3_1313_728 = lever[4] & lever[25];
assign xor_1282_774 = gate3_1214_728 ^ gate3_1304_728;
assign gate3_1304_728 = lever[5] & lever[24];
assign gate3_1214_728 = lever[23] & lever[6];
assign gate3_1279_774 = gate3_1214_728 & gate3_1304_728;
assign gate3_16_1054 = not_1140_858 | not_17_1053;
assign not_17_1053 = ~gate3_599_983;
assign xor_23_1453 = not_23_1395 ^ gate3_17_1430;
assign gate3_17_1430 = gate3_7_1366 | not_18_1429;
assign not_18_1429 = ~gate3_17_1394;
assign gate3_17_1394 = not_18_1234 | not_18_1393;
assign not_18_1393 = ~not_20_1367;
assign not_20_1367 = ~xor_20_1366;
assign xor_20_1366 = gate3_7_1330 ^ not_22_1280;
assign not_22_1280 = ~xor_22_1279;
assign xor_22_1279 = not_22_1234 ^ xor_24_1108;
assign gate3_7_1330 = gate3_3_1233 & gate3_1_1279;
assign gate3_1_1279 = not_2_1278 | xor_1_1108;
assign xor_1_1108 = gate3_1_983 ^ xor_7_1054;
assign not_2_1278 = ~not_6_1234;
assign not_6_1234 = ~xor_6_1233;
assign xor_6_1233 = gate3_3_1182 ^ xor_12_1108;
assign xor_12_1108 = not_3_858 ^ xor_13_1054;
assign gate3_3_1182 = gate3_7_1108 & gate3_10_1054;
assign gate3_10_1054 = not_1134_858 | not_11_1053;
assign not_11_1053 = ~gate3_596_983;
assign gate3_596_983 = gate3_1104_857 | gate3_1264_774;
assign gate3_1264_774 = gate3_1202_728 & gate3_1277_728;
assign gate3_1277_728 = lever[21] & lever[7];
assign gate3_1202_728 = lever[20] & lever[8];
assign gate3_1104_857 = xor_1267_774 & gate3_1307_728;
assign gate3_1307_728 = lever[22] & lever[6];
assign xor_1267_774 = gate3_1202_728 ^ gate3_1277_728;
assign not_1134_858 = ~xor_1134_857;
assign xor_1134_857 = gate3_1205_728 ^ xor_1174_774;
assign gate3_7_1108 = not_1128_858 | xor_728_1054;
assign xor_728_1054 = gate3_596_983 ^ not_1134_858;
assign not_1128_858 = ~xor_1128_857;
assign xor_1128_857 = gate3_1313_728 ^ xor_1282_774;
assign gate3_3_1233 = not_4_1232 | gate3_3_1182;
assign not_4_1232 = ~xor_12_1108;
assign not_18_1234 = ~xor_18_1233;
assign xor_18_1233 = not_5_984 ^ gate3_7_1182;
assign gate3_7_1366 = not_22_1280 & not_8_1365;
assign not_8_1365 = ~gate3_7_1330;
assign not_23_1395 = ~xor_23_1394;
assign xor_23_1394 = xor_25_1279 ^ xor_23_1366;
assign gate3_20_1453 = not_23_1395 | not_21_1452;
assign not_21_1452 = ~gate3_17_1430;
assign xor_45_1528 = gate3_36_1503 ^ not_47_1479;
assign gate3_17_1555 = gate3_12_1528 & not_42_1529;
assign not_42_1529 = ~xor_42_1528;
assign xor_42_1528 = xor_44_1478 ^ gate3_33_1503;
assign gate3_12_1528 = xor_25_1478 & gate3_7_1503;
assign gate3_7_1503 = not_8_1502 | gate3_10_1453;
assign gate3_10_1453 = gate3_5_1430 & not_20_1395;
assign not_20_1395 = ~xor_20_1394;
assign xor_20_1394 = not_18_1234 ^ not_20_1367;
assign gate3_5_1430 = gate3_1_1366 | not_6_1429;
assign not_6_1429 = ~gate3_3_1394;
assign gate3_3_1394 = not_4_1393 | xor_9_1233;
assign xor_9_1233 = gate3_448_1182 ^ xor_1285_774;
assign xor_1285_774 = gate3_1193_728 ^ gate3_1226_728;
assign gate3_1226_728 = lever[0] & lever[30];
assign gate3_1193_728 = lever[29] & lever[1];
assign gate3_448_1182 = gate3_722_1054 & gate3_760_1108;
assign gate3_760_1108 = xor_725_1054 | not_761_1107;
assign not_761_1107 = ~gate3_587_983;
assign gate3_587_983 = gate3_1246_774 | gate3_1086_857;
assign gate3_1086_857 = gate3_1289_728 & xor_1252_774;
assign xor_1252_774 = gate3_1286_728 ^ gate3_1292_728;
assign gate3_1292_728 = lever[2] & lever[26];
assign gate3_1286_728 = lever[1] & lever[27];
assign gate3_1289_728 = lever[0] & lever[28];
assign gate3_1246_774 = gate3_1286_728 & gate3_1292_728;
assign xor_725_1054 = not_1116_858 ^ gate3_590_983;
assign gate3_590_983 = gate3_1255_774 | gate3_1092_857;
assign gate3_1092_857 = gate3_1298_728 & xor_1258_774;
assign xor_1258_774 = gate3_1301_728 ^ gate3_1268_728;
assign gate3_1268_728 = lever[4] & lever[24];
assign gate3_1301_728 = lever[23] & lever[5];
assign gate3_1298_728 = lever[3] & lever[25];
assign gate3_1255_774 = gate3_1268_728 & gate3_1301_728;
assign not_1116_858 = ~xor_1116_857;
assign xor_1116_857 = gate3_1310_728 ^ xor_1276_774;
assign gate3_722_1054 = not_723_1053 | not_1116_858;
assign not_723_1053 = ~gate3_590_983;
assign not_4_1393 = ~xor_4_1366;
assign xor_4_1366 = not_5_1280 ^ gate3_1_1330;
assign gate3_1_1330 = gate3_512_1233 | not_2_1329;
assign not_2_1329 = ~gate3_556_1279;
assign gate3_556_1279 = xor_763_1108 | not_557_1278;
assign not_557_1278 = ~not_515_1234;
assign not_515_1234 = ~xor_515_1233;
assign xor_515_1233 = gate3_439_1182 ^ xor_766_1108;
assign xor_766_1108 = not_1128_858 ^ xor_728_1054;
assign gate3_439_1182 = gate3_754_1108 & gate3_716_1054;
assign gate3_716_1054 = not_1107_858 | not_717_1053;
assign not_717_1053 = ~gate3_584_983;
assign gate3_584_983 = gate3_1231_774 | gate3_1077_857;
assign gate3_1077_857 = xor_1234_774 & gate3_1271_728;
assign gate3_1271_728 = lever[22] & lever[5];
assign xor_1234_774 = gate3_1274_728 ^ gate3_1247_728;
assign gate3_1247_728 = lever[21] & lever[6];
assign gate3_1274_728 = lever[20] & lever[7];
assign gate3_1231_774 = gate3_1247_728 & gate3_1274_728;
assign not_1107_858 = ~xor_1107_857;
assign xor_1107_857 = gate3_1307_728 ^ xor_1267_774;
assign gate3_754_1108 = xor_719_1054 | not_1098_858;
assign not_1098_858 = ~xor_1098_857;
assign xor_1098_857 = gate3_1298_728 ^ xor_1258_774;
assign xor_719_1054 = not_1107_858 ^ gate3_584_983;
assign xor_763_1108 = gate3_587_983 ^ xor_725_1054;
assign gate3_512_1233 = not_513_1232 & xor_766_1108;
assign not_513_1232 = ~gate3_439_1182;
assign not_5_1280 = ~xor_5_1279;
assign xor_5_1279 = xor_1_1108 ^ not_6_1234;
assign gate3_1_1366 = gate3_1_1330 & not_5_1280;
assign not_8_1502 = ~gate3_15_1478;
assign gate3_15_1478 = not_17_1454 | gate3_28_1233;
assign gate3_28_1233 = gate3_448_1182 | not_29_1232;
assign not_29_1232 = ~xor_1285_774;
assign not_17_1454 = ~xor_17_1453;
assign xor_17_1453 = gate3_5_1430 ^ not_20_1395;
assign xor_25_1478 = gate3_15_1233 ^ xor_23_1453;
assign xor_24_1576 = gate3_51_1528 ^ not_37_1556;
assign gate3_20_1602 = gate3_28_1555 & xor_24_1576;
assign gate3_28_1555 = gate3_38_1528 & xor_45_1528;
assign not_2_1727 = ~gate3_1_1720;
assign gate3_1_1720 = gate3_1_1714 | gate3_19_1628;
assign gate3_19_1628 = not_24_1603 | gate3_27_1602;
assign gate3_27_1602 = gate3_30_1576 | not_28_1601;
assign not_28_1601 = ~gate3_37_1576;
assign gate3_37_1576 = gate3_17_1555 | not_38_1575;
assign not_38_1575 = ~not_40_1556;
assign not_24_1603 = ~xor_24_1602;
assign xor_24_1602 = xor_24_1576 ^ gate3_28_1555;
assign gate3_1_1714 = not_2_1713 & gate3_6_1654;
assign gate3_6_1654 = gate3_10_1602 & gate3_6_1628;
assign gate3_6_1628 = gate3_1_1602 | not_22_1556;
assign not_22_1556 = ~xor_22_1555;
assign xor_22_1555 = gate3_12_1528 ^ not_42_1529;
assign gate3_1_1602 = gate3_4_1555 | not_6_1577;
assign not_6_1577 = ~xor_6_1576;
assign xor_6_1576 = gate3_1_1555 ^ not_15_1529;
assign not_15_1529 = ~xor_15_1528;
assign xor_15_1528 = gate3_7_1503 ^ xor_25_1478;
assign gate3_1_1555 = not_4_1528 | not_2_1554;
assign not_2_1554 = ~xor_18_1478;
assign xor_18_1478 = gate3_28_1233 ^ not_17_1454;
assign not_4_1528 = ~gate3_4_1503;
assign gate3_4_1503 = gate3_1_1453 | not_5_1502;
assign not_5_1502 = ~gate3_3_1478;
assign gate3_3_1478 = not_4_1454 | gate3_12_1233;
assign gate3_12_1233 = not_13_1232 | gate3_436_1182;
assign gate3_436_1182 = not_437_1181 & gate3_707_1054;
assign gate3_707_1054 = not_1089_858 | not_708_1053;
assign not_708_1053 = ~gate3_581_983;
assign gate3_581_983 = gate3_1219_774 | gate3_1068_857;
assign gate3_1068_857 = gate3_1262_728 & xor_1225_774;
assign xor_1225_774 = gate3_1259_728 ^ gate3_1265_728;
assign gate3_1265_728 = lever[23] & lever[4];
assign gate3_1259_728 = lever[24] & lever[3];
assign gate3_1262_728 = lever[2] & lever[25];
assign gate3_1219_774 = gate3_1259_728 & gate3_1265_728;
assign not_1089_858 = ~xor_1089_857;
assign xor_1089_857 = gate3_1289_728 ^ xor_1252_774;
assign not_437_1181 = ~gate3_745_1108;
assign gate3_745_1108 = gate3_1237_774 & not_746_1107;
assign not_746_1107 = ~xor_710_1054;
assign xor_710_1054 = not_1089_858 ^ gate3_581_983;
assign gate3_1237_774 = gate3_1286_728 & gate3_28_728;
assign gate3_28_728 = lever[0] & lever[26];
assign not_13_1232 = ~gate3_1229_728;
assign not_4_1454 = ~xor_4_1453;
assign xor_4_1453 = gate3_2_1430 ^ not_9_1395;
assign not_9_1395 = ~xor_9_1394;
assign xor_9_1394 = xor_9_1233 ^ xor_4_1366;
assign gate3_2_1430 = gate3_389_1366 | gate3_406_1394;
assign gate3_406_1394 = not_509_1234 & not_407_1393;
assign not_407_1393 = ~not_393_1367;
assign not_393_1367 = ~xor_393_1366;
assign xor_393_1366 = gate3_352_1330 ^ not_559_1280;
assign not_559_1280 = ~xor_559_1279;
assign xor_559_1279 = xor_763_1108 ^ not_515_1234;
assign gate3_352_1330 = gate3_503_1233 | not_353_1329;
assign not_353_1329 = ~gate3_550_1279;
assign gate3_550_1279 = not_551_1278 | xor_748_1108;
assign xor_748_1108 = gate3_1237_774 ^ xor_710_1054;
assign not_551_1278 = ~not_506_1234;
assign not_506_1234 = ~xor_506_1233;
assign xor_506_1233 = xor_757_1108 ^ gate3_432_1182;
assign gate3_432_1182 = gate3_700_1054 & gate3_739_1108;
assign gate3_739_1108 = xor_704_1054 | not_1074_858;
assign not_1074_858 = ~xor_1074_857;
assign xor_1074_857 = gate3_1262_728 ^ xor_1225_774;
assign xor_704_1054 = not_1080_858 ^ gate3_575_983;
assign gate3_575_983 = gate3_1201_774 | gate3_1056_857;
assign gate3_1056_857 = gate3_1241_728 & xor_1210_774;
assign xor_1210_774 = gate3_1238_728 ^ gate3_1244_728;
assign gate3_1244_728 = lever[20] & lever[6];
assign gate3_1238_728 = lever[21] & lever[5];
assign gate3_1241_728 = lever[22] & lever[4];
assign gate3_1201_774 = gate3_1238_728 & gate3_1244_728;
assign not_1080_858 = ~xor_1080_857;
assign xor_1080_857 = gate3_1271_728 ^ xor_1234_774;
assign gate3_700_1054 = not_1080_858 | not_701_1053;
assign not_701_1053 = ~gate3_575_983;
assign xor_757_1108 = not_1098_858 ^ xor_719_1054;
assign gate3_503_1233 = not_504_1232 & xor_757_1108;
assign not_504_1232 = ~gate3_432_1182;
assign not_509_1234 = ~xor_509_1233;
assign xor_509_1233 = gate3_1229_728 ^ gate3_436_1182;
assign gate3_389_1366 = gate3_352_1330 & not_559_1280;
assign gate3_1_1453 = gate3_2_1430 & not_9_1395;
assign gate3_4_1555 = gate3_1_1503 | not_6_1529;
assign not_6_1529 = ~xor_6_1528;
assign xor_6_1528 = gate3_4_1503 ^ xor_18_1478;
assign gate3_1_1503 = gate3_7_1453 | not_12_1479;
assign not_12_1479 = ~xor_12_1478;
assign xor_12_1478 = gate3_12_1233 ^ not_4_1454;
assign gate3_7_1453 = xor_35_1394 | not_8_1452;
assign not_8_1452 = ~gate3_30_1430;
assign gate3_30_1430 = gate3_386_1366 | gate3_403_1394;
assign gate3_403_1394 = gate3_49_1054 & not_404_1393;
assign not_404_1393 = ~not_36_1367;
assign not_36_1367 = ~xor_36_1366;
assign xor_36_1366 = gate3_349_1330 ^ not_553_1280;
assign not_553_1280 = ~xor_553_1279;
assign xor_553_1279 = xor_748_1108 ^ not_506_1234;
assign gate3_349_1330 = gate3_547_1279 | gate3_500_1233;
assign gate3_500_1233 = xor_742_1108 & not_501_1232;
assign not_501_1232 = ~gate3_429_1182;
assign gate3_429_1182 = gate3_736_1108 & gate3_697_1054;
assign gate3_697_1054 = not_1059_858 | not_698_1053;
assign not_698_1053 = ~gate3_569_983;
assign gate3_569_983 = gate3_1050_857 | gate3_1198_774;
assign gate3_1198_774 = gate3_1232_728 & gate3_1235_728;
assign gate3_1235_728 = lever[20] & lever[5];
assign gate3_1232_728 = lever[21] & lever[4];
assign gate3_1050_857 = gate3_13_728 & xor_7_774;
assign xor_7_774 = gate3_1232_728 ^ gate3_1235_728;
assign gate3_13_728 = lever[22] & lever[3];
assign not_1059_858 = ~xor_1059_857;
assign xor_1059_857 = gate3_1241_728 ^ xor_1210_774;
assign gate3_736_1108 = not_30_858 | xor_28_1054;
assign xor_28_1054 = gate3_569_983 ^ not_1059_858;
assign not_30_858 = ~xor_30_857;
assign xor_30_857 = gate3_1250_728 ^ xor_1216_774;
assign xor_1216_774 = gate3_1253_728 ^ gate3_1256_728;
assign gate3_1256_728 = lever[3] & lever[23];
assign gate3_1253_728 = lever[2] & lever[24];
assign gate3_1250_728 = lever[1] & lever[25];
assign xor_742_1108 = not_1074_858 ^ xor_704_1054;
assign gate3_547_1279 = xor_45_1054 & not_43_1234;
assign not_43_1234 = ~xor_43_1233;
assign xor_43_1233 = xor_742_1108 ^ gate3_429_1182;
assign xor_45_1054 = xor_1243_774 ^ gate3_578_983;
assign gate3_578_983 = gate3_1213_774 | gate3_1065_857;
assign gate3_1065_857 = gate3_1250_728 & xor_1216_774;
assign gate3_1213_774 = gate3_1253_728 & gate3_1256_728;
assign xor_1243_774 = gate3_1280_728 ^ gate3_1283_728;
assign gate3_1283_728 = lever[0] & lever[27];
assign gate3_1280_728 = lever[1] & lever[26];
assign gate3_49_1054 = xor_1243_774 & gate3_578_983;
assign gate3_386_1366 = gate3_349_1330 & not_553_1280;
assign xor_35_1394 = not_509_1234 ^ not_393_1367;
assign gate3_10_1602 = gate3_1_1576 | not_22_1556;
assign gate3_1_1576 = gate3_1_1555 | not_15_1529;
assign not_2_1713 = ~gate3_1_1706;
assign gate3_1_1706 = gate3_1_1693 & xor_17_1602;
assign xor_17_1602 = gate3_1_1576 ^ not_22_1556;
assign gate3_1_1693 = gate3_1_1679 & xor_4_1602;
assign xor_4_1602 = gate3_4_1555 ^ not_6_1577;
assign gate3_1_1679 = gate3_12_1576 | gate3_1_1654;
assign gate3_1_1654 = xor_15_1576 & gate3_1_1628;
assign gate3_1_1628 = gate3_7_1602 | gate3_35_1528;
assign gate3_35_1528 = xor_10_1503 & not_36_1527;
assign not_36_1527 = ~gate3_13_1503;
assign gate3_13_1503 = not_14_1502 | gate3_31_1478;
assign gate3_31_1478 = gate3_37_1430 | xor_33_1453;
assign xor_33_1453 = gate3_25_1430 ^ xor_32_1394;
assign xor_32_1394 = gate3_49_1054 ^ not_36_1367;
assign gate3_25_1430 = gate3_30_1366 | gate3_26_1394;
assign gate3_26_1394 = gate3_38_1054 & not_27_1393;
assign not_27_1393 = ~not_33_1367;
assign not_33_1367 = ~xor_33_1366;
assign xor_33_1366 = xor_36_1279 ^ gate3_30_1330;
assign gate3_30_1330 = gate3_31_1233 | gate3_33_1279;
assign gate3_33_1279 = xor_41_1054 & not_35_1234;
assign not_35_1234 = ~xor_35_1233;
assign xor_35_1233 = gate3_10_1182 ^ xor_30_1108;
assign xor_30_1108 = not_30_858 ^ xor_28_1054;
assign gate3_10_1182 = gate3_19_1054 & gate3_27_1108;
assign gate3_27_1108 = not_26_858 | xor_22_1054;
assign xor_22_1054 = gate3_8_983 ^ not_15_858;
assign not_15_858 = ~xor_15_857;
assign xor_15_857 = gate3_13_728 ^ xor_7_774;
assign gate3_8_983 = gate3_1_774 | gate3_12_857;
assign gate3_12_857 = gate3_10_728 & xor_4_774;
assign xor_4_774 = gate3_1_728 ^ gate3_7_728;
assign gate3_7_728 = lever[4] & lever[20];
assign gate3_1_728 = lever[21] & lever[3];
assign gate3_10_728 = lever[2] & lever[22];
assign gate3_1_774 = gate3_1_728 & gate3_7_728;
assign not_26_858 = ~xor_26_857;
assign xor_26_857 = gate3_16_728 ^ xor_21_774;
assign xor_21_774 = gate3_25_728 ^ gate3_19_728;
assign gate3_19_728 = lever[24] & lever[1];
assign gate3_25_728 = lever[23] & lever[2];
assign gate3_16_728 = lever[0] & lever[25];
assign gate3_19_1054 = not_20_1053 | not_15_858;
assign not_20_1053 = ~gate3_8_983;
assign xor_41_1054 = gate3_11_983 ^ gate3_28_728;
assign gate3_11_983 = gate3_18_774 | gate3_20_857;
assign gate3_20_857 = gate3_16_728 & xor_21_774;
assign gate3_18_774 = gate3_19_728 & gate3_25_728;
assign gate3_31_1233 = xor_30_1108 & not_32_1232;
assign not_32_1232 = ~gate3_10_1182;
assign xor_36_1279 = xor_45_1054 ^ not_43_1234;
assign gate3_38_1054 = gate3_11_983 & gate3_28_728;
assign gate3_30_1366 = gate3_30_1330 & xor_36_1279;
assign gate3_37_1430 = xor_38_1394 | not_42_1394;
assign not_42_1394 = ~gate3_42_1366;
assign gate3_42_1366 = gate3_33_1330 & not_43_1365;
assign not_43_1365 = ~not_43_1280;
assign not_43_1280 = ~xor_43_1279;
assign xor_43_1279 = xor_41_1054 ^ not_35_1234;
assign gate3_33_1330 = gate3_47_1233 | gate3_40_1279;
assign gate3_40_1279 = not_51_1234 & gate3_33_774;
assign gate3_33_774 = gate3_19_728 & gate3_47_728;
assign gate3_47_728 = lever[0] & lever[23];
assign not_51_1234 = ~xor_51_1233;
assign xor_51_1233 = gate3_14_1182 ^ xor_43_1108;
assign xor_43_1108 = not_26_858 ^ xor_22_1054;
assign gate3_14_1182 = gate3_52_1054 & gate3_35_1108;
assign gate3_35_1108 = not_36_775 | xor_55_1054;
assign xor_55_1054 = gate3_17_983 ^ not_41_858;
assign not_41_858 = ~xor_41_857;
assign xor_41_857 = gate3_10_728 ^ xor_4_774;
assign gate3_17_983 = gate3_24_774 | gate3_38_857;
assign gate3_38_857 = xor_30_774 & gate3_41_728;
assign gate3_41_728 = lever[1] & lever[22];
assign xor_30_774 = gate3_31_728 ^ gate3_4_728;
assign gate3_4_728 = lever[20] & lever[3];
assign gate3_31_728 = lever[21] & lever[2];
assign gate3_24_774 = gate3_1_728 & gate3_34_728;
assign gate3_34_728 = lever[20] & lever[2];
assign not_36_775 = ~xor_36_774;
assign xor_36_774 = gate3_22_728 ^ gate3_44_728;
assign gate3_44_728 = lever[24] & lever[0];
assign gate3_22_728 = lever[1] & lever[23];
assign gate3_52_1054 = not_53_1053 | not_41_858;
assign not_53_1053 = ~gate3_17_983;
assign gate3_47_1233 = xor_43_1108 & not_48_1232;
assign not_48_1232 = ~gate3_14_1182;
assign xor_38_1394 = gate3_38_1054 ^ not_33_1367;
assign not_14_1502 = ~xor_34_1478;
assign xor_34_1478 = gate3_26_1453 ^ xor_30_1453;
assign xor_30_1453 = xor_35_1394 ^ gate3_30_1430;
assign gate3_26_1453 = xor_32_1394 | not_27_1452;
assign not_27_1452 = ~gate3_25_1430;
assign xor_10_1503 = gate3_7_1453 ^ not_12_1479;
assign gate3_7_1602 = gate3_18_1576 & not_10_1556;
assign not_10_1556 = ~xor_10_1555;
assign xor_10_1555 = xor_10_1503 ^ gate3_23_1528;
assign gate3_23_1528 = gate3_13_1503 & gate3_28_1478;
assign gate3_28_1478 = xor_30_1453 | gate3_26_1453;
assign gate3_18_1576 = gate3_26_1528 | gate3_13_1555;
assign gate3_13_1555 = gate3_29_1528 & gate3_32_1528;
assign gate3_32_1528 = gate3_23_1503 & xor_30_1503;
assign xor_30_1503 = gate3_42_1453 ^ xor_37_1478;
assign xor_37_1478 = gate3_37_1430 ^ xor_33_1453;
assign gate3_42_1453 = not_44_1430 & not_43_1452;
assign not_43_1452 = ~not_40_1431;
assign not_40_1431 = ~xor_40_1430;
assign xor_40_1430 = not_42_1394 ^ xor_38_1394;
assign not_44_1430 = ~gate3_44_1394;
assign gate3_44_1394 = xor_45_1366 | gate3_40_1330;
assign gate3_40_1330 = not_51_1280 | gate3_54_1233;
assign gate3_54_1233 = gate3_17_1182 | not_55_1232;
assign not_55_1232 = ~xor_54_1108;
assign xor_54_1108 = not_36_775 ^ xor_55_1054;
assign gate3_17_1182 = not_18_1181 & gate3_87_1054;
assign gate3_87_1054 = not_88_1053 | not_52_858;
assign not_52_858 = ~xor_52_857;
assign xor_52_857 = gate3_41_728 ^ xor_30_774;
assign not_88_1053 = ~gate3_20_983;
assign gate3_20_983 = gate3_43_774 | gate3_45_857;
assign gate3_45_857 = gate3_53_728 & xor_88_774;
assign xor_88_774 = gate3_34_728 ^ gate3_50_728;
assign gate3_50_728 = lever[1] & lever[21];
assign gate3_53_728 = lever[0] & lever[22];
assign gate3_43_774 = gate3_50_728 & gate3_34_728;
assign not_18_1181 = ~gate3_47_1108;
assign gate3_47_1108 = gate3_47_728 & not_48_1107;
assign not_48_1107 = ~xor_95_1054;
assign xor_95_1054 = gate3_20_983 ^ not_52_858;
assign not_51_1280 = ~xor_51_1279;
assign xor_51_1279 = gate3_33_774 ^ not_51_1234;
assign xor_45_1366 = not_43_1280 ^ gate3_33_1330;
assign gate3_23_1503 = gate3_56_1366 & gate3_40_1478;
assign gate3_40_1478 = not_40_1453 & xor_47_1394;
assign xor_47_1394 = xor_45_1366 ^ gate3_40_1330;
assign not_40_1453 = ~not_40_1431;
assign gate3_56_1366 = gate3_20_1182 & not_57_1365;
assign not_57_1365 = ~gate3_45_1330;
assign gate3_45_1330 = not_51_1280 | not_46_1329;
assign not_46_1329 = ~not_85_1234;
assign not_85_1234 = ~xor_85_1233;
assign xor_85_1233 = gate3_17_1182 ^ xor_54_1108;
assign gate3_20_1182 = not_57_1109 & gate3_98_1054;
assign gate3_98_1054 = gate3_23_983 & gate3_56_728;
assign gate3_56_728 = lever[20] & lever[0];
assign gate3_23_983 = gate3_50_728 & not_24_982;
assign not_24_982 = ~not_85_858;
assign not_85_858 = ~xor_85_857;
assign xor_85_857 = gate3_53_728 ^ xor_88_774;
assign not_57_1109 = ~xor_57_1108;
assign xor_57_1108 = gate3_47_728 ^ xor_95_1054;
assign gate3_29_1528 = not_20_1504 | gate3_16_1503;
assign gate3_16_1503 = gate3_42_1453 & xor_37_1478;
assign not_20_1504 = ~xor_20_1503;
assign xor_20_1503 = gate3_31_1478 ^ xor_34_1478;
assign gate3_26_1528 = gate3_16_1503 & not_20_1504;
assign xor_15_1576 = xor_7_1555 ^ gate3_20_1528;
assign gate3_20_1528 = not_28_1503 & xor_10_1503;
assign not_28_1503 = ~gate3_28_1478;
assign xor_7_1555 = not_6_1529 ^ gate3_1_1503;
assign gate3_12_1576 = gate3_20_1528 & xor_7_1555;
assign gate3_62_1628 = not_43_1577 & not_63_1627;
assign not_63_1627 = ~gate3_54_1602;
assign gate3_92_1628 = xor_84_1602 | xor_90_1602;
assign xor_90_1602 = gate3_66_1576 ^ not_77_1556;
assign gate3_1_1915 = gate3_1_1908 | xor_69_1576;
assign gate3_7_1915 = gate3_6_1908 & not_8_1914;
assign not_8_1914 = ~gate3_4_1901;
assign gate3_4_1901 = xor_90_1602 & gate3_1_1892;
assign gate3_6_1908 = gate3_7_1901 & gate3_10_1901;
assign gate3_10_1901 = gate3_4_1892 & not_11_1900;
assign not_11_1900 = ~gate3_7_1892;
assign gate3_7_1892 = gate3_9_1885 | not_8_1891;
assign not_8_1891 = ~gate3_12_1885;
assign gate3_12_1885 = gate3_1_1876 | gate3_129_1654;
assign gate3_129_1654 = gate3_77_1628 & not_130_1653;
assign not_130_1653 = ~gate3_87_1628;
assign gate3_9_1885 = gate3_1_1876 & gate3_117_1654;
assign gate3_117_1654 = gate3_77_1628 & gate3_84_1628;
assign gate3_4_1892 = not_5_1891 & gate3_6_1885;
assign gate3_6_1885 = gate3_10_1876 & gate3_7_1876;
assign gate3_7_1876 = not_8_1875 | gate3_75_1654;
assign gate3_75_1654 = gate3_62_1628 | not_76_1653;
assign not_76_1653 = ~gate3_59_1628;
assign not_8_1875 = ~gate3_6_1866;
assign gate3_6_1866 = gate3_111_1679 & gate3_1_1857;
assign gate3_10_1876 = gate3_9_1866 & not_4_1858;
assign not_4_1858 = ~xor_4_1857;
assign xor_4_1857 = xor_108_1679 ^ gate3_1_1849;
assign gate3_9_1866 = gate3_10_1857 & not_10_1865;
assign not_10_1865 = ~gate3_7_1857;
assign gate3_7_1857 = gate3_6_1849 & gate3_84_1693;
assign gate3_84_1693 = xor_86_1679 | not_85_1692;
assign not_85_1692 = ~gate3_105_1679;
assign gate3_6_1849 = not_7_1848 | gate3_6_1841;
assign gate3_6_1841 = gate3_1_1834 & gate3_94_1679;
assign not_7_1848 = ~gate3_9_1841;
assign gate3_9_1841 = not_10_1840 | gate3_1_1834;
assign not_10_1840 = ~gate3_16_1706;
assign gate3_10_1857 = gate3_9_1849 & gate3_4_1834;
assign gate3_4_1834 = not_9_1828 & gate3_4_1819;
assign gate3_4_1819 = not_4_1814 & gate3_9_1800;
assign gate3_9_1800 = not_10_1799 & gate3_12_1793;
assign gate3_12_1793 = gate3_13_1785 & not_13_1792;
assign not_13_1792 = ~gate3_9_1778;
assign gate3_9_1778 = not_14_1655 & gate3_1_1770;
assign gate3_13_1785 = gate3_1_1778 & gate3_13_1778;
assign gate3_13_1778 = gate3_18_1764 & gate3_9_1770;
assign gate3_9_1770 = gate3_20_1743 & gate3_22_1764;
assign gate3_22_1764 = gate3_22_1756 & gate3_18_1728;
assign gate3_18_1728 = not_19_1727 | gate3_30_1576;
assign not_19_1727 = ~gate3_18_1720;
assign gate3_18_1720 = gate3_1_1714 & gate3_103_1628;
assign gate3_103_1628 = not_24_1603 | gate3_37_1576;
assign gate3_22_1756 = gate3_22_1749 & gate3_47_1714;
assign gate3_47_1714 = gate3_48_1706 & not_48_1713;
assign not_48_1713 = ~gate3_88_1693;
assign gate3_88_1693 = xor_43_1679 & gate3_46_1679;
assign gate3_48_1706 = gate3_4_1693 & gate3_119_1693;
assign gate3_119_1693 = gate3_131_1679 & not_120_1692;
assign not_120_1692 = ~gate3_84_1654;
assign gate3_84_1654 = xor_41_1628 & not_85_1653;
assign not_85_1653 = ~gate3_37_1628;
assign gate3_131_1679 = not_94_1655 & gate3_87_1654;
assign gate3_87_1654 = gate3_98_1602 | gate3_106_1628;
assign gate3_106_1628 = gate3_104_1602 | not_107_1627;
assign not_107_1627 = ~gate3_79_1576;
assign gate3_79_1576 = not_80_1575 | not_113_1529;
assign not_80_1575 = ~gate3_84_1555;
assign gate3_104_1602 = xor_96_1576 | gate3_99_1576;
assign gate3_99_1576 = xor_131_1528 & gate3_92_1555;
assign gate3_92_1555 = gate3_89_1503 | gate3_118_1528;
assign gate3_118_1528 = not_92_1504 & gate3_104_728;
assign gate3_104_728 = lever[15] & lever[39];
assign not_92_1504 = ~xor_92_1503;
assign xor_92_1503 = gate3_95_1478 ^ not_121_1454;
assign not_121_1454 = ~xor_121_1453;
assign xor_121_1453 = xor_127_1366 ^ gate3_116_1430;
assign gate3_116_1430 = gate3_116_1366 & not_117_1429;
assign not_117_1429 = ~gate3_111_1394;
assign gate3_111_1394 = not_112_1393 & gate3_101_728;
assign not_112_1393 = ~xor_121_1366;
assign gate3_116_1366 = not_111_1280 | not_117_1365;
assign not_117_1365 = ~gate3_95_1330;
assign xor_127_1366 = not_133_1234 ^ gate3_98_1330;
assign gate3_98_1330 = gate3_121_1233 | gate3_106_1279;
assign gate3_106_1279 = gate3_83_728 & not_124_1234;
assign gate3_121_1233 = gate3_51_1182 & not_122_1232;
assign not_122_1232 = ~xor_115_1054;
assign not_133_1234 = ~xor_133_1233;
assign xor_133_1233 = gate3_107_728 ^ not_85_1183;
assign not_85_1183 = ~xor_85_1182;
assign xor_85_1182 = gate3_111_1108 ^ xor_141_1054;
assign xor_141_1054 = not_117_858 ^ gate3_54_983;
assign gate3_54_983 = gate3_94_774 | gate3_96_857;
assign gate3_96_857 = xor_97_774 & gate3_86_728;
assign gate3_94_774 = gate3_95_728 & gate3_92_728;
assign gate3_92_728 = lever[18] & lever[36];
assign not_117_858 = ~xor_117_857;
assign xor_117_857 = xor_124_774 ^ gate3_110_728;
assign gate3_110_728 = lever[17] & lever[37];
assign xor_124_774 = gate3_113_728 ^ gate3_92_728;
assign gate3_113_728 = lever[19] & lever[35];
assign gate3_111_1108 = gate3_112_1054 | gate3_43_983;
assign gate3_43_983 = gate3_112_774 & not_44_982;
assign not_44_982 = ~not_99_858;
assign gate3_112_1054 = gate3_38_983 & not_113_1053;
assign not_113_1053 = ~xor_49_983;
assign gate3_107_728 = lever[16] & lever[38];
assign gate3_95_1478 = gate3_106_1453 | not_96_1477;
assign not_96_1477 = ~gate3_111_1453;
assign gate3_111_1453 = not_112_1452 | gate3_106_1394;
assign not_112_1452 = ~xor_111_1430;
assign gate3_106_1453 = not_121_1430 & not_107_1452;
assign not_107_1452 = ~xor_114_1394;
assign not_121_1430 = ~gate3_121_1394;
assign gate3_89_1503 = gate3_95_1478 & not_90_1502;
assign not_90_1502 = ~not_121_1454;
assign xor_131_1528 = not_95_1504 ^ gate3_119_728;
assign gate3_119_728 = lever[16] & lever[39];
assign not_95_1504 = ~xor_95_1503;
assign xor_95_1503 = gate3_99_1478 ^ xor_109_1330;
assign xor_109_1330 = xor_95_1182 ^ gate3_123_1279;
assign gate3_123_1279 = gate3_129_1233 | gate3_56_1182;
assign gate3_56_1182 = gate3_111_1108 & not_57_1181;
assign not_57_1181 = ~xor_141_1054;
assign gate3_129_1233 = gate3_107_728 & not_85_1183;
assign xor_95_1182 = gate3_122_728 ^ xor_124_1108;
assign xor_124_1108 = gate3_124_1054 ^ not_148_1055;
assign not_148_1055 = ~xor_148_1054;
assign xor_148_1054 = gate3_87_983 ^ xor_148_774;
assign xor_148_774 = gate3_125_728 ^ gate3_116_728;
assign gate3_116_728 = lever[36] & lever[19];
assign gate3_125_728 = lever[18] & lever[37];
assign gate3_87_983 = gate3_115_774 | gate3_109_857;
assign gate3_109_857 = gate3_110_728 & xor_124_774;
assign gate3_115_774 = gate3_89_728 & gate3_116_728;
assign gate3_124_1054 = not_125_1053 & gate3_54_983;
assign not_125_1053 = ~not_117_858;
assign gate3_122_728 = lever[17] & lever[38];
assign gate3_99_1478 = not_124_1394 | gate3_117_1453;
assign gate3_117_1453 = not_118_1452 & not_127_1394;
assign not_127_1394 = ~xor_127_1366;
assign not_118_1452 = ~gate3_116_1430;
assign not_124_1394 = ~gate3_124_1366;
assign gate3_124_1366 = not_133_1234 | not_125_1365;
assign not_125_1365 = ~gate3_98_1330;
assign xor_96_1576 = gate3_99_1555 ^ not_111_1479;
assign not_111_1479 = ~xor_111_1478;
assign xor_111_1478 = gate3_131_728 ^ xor_133_1453;
assign xor_133_1453 = xor_139_1366 ^ gate3_133_1430;
assign gate3_133_1430 = not_124_1394 & not_134_1429;
assign not_134_1429 = ~xor_109_1330;
assign xor_139_1366 = gate3_106_1330 ^ xor_135_1279;
assign xor_135_1279 = gate3_139_1233 ^ xor_112_1182;
assign xor_112_1182 = not_139_1109 ^ gate3_134_728;
assign gate3_134_728 = lever[18] & lever[38];
assign not_139_1109 = ~xor_139_1108;
assign xor_139_1108 = gate3_151_774 ^ gate3_145_1054;
assign gate3_145_1054 = xor_148_774 & gate3_87_983;
assign gate3_151_774 = gate3_128_728 & not_152_773;
assign not_152_773 = ~gate3_92_728;
assign gate3_128_728 = lever[37] & lever[19];
assign gate3_139_1233 = gate3_117_1108 | gate3_88_1182;
assign gate3_88_1182 = not_89_1181 & gate3_122_728;
assign not_89_1181 = ~xor_124_1108;
assign gate3_117_1108 = gate3_124_1054 & not_118_1107;
assign not_118_1107 = ~not_148_1055;
assign gate3_106_1330 = xor_95_1182 | not_107_1329;
assign not_107_1329 = ~gate3_123_1279;
assign gate3_131_728 = lever[17] & lever[39];
assign gate3_99_1555 = gate3_102_1478 | gate3_125_1528;
assign gate3_125_1528 = not_95_1504 & gate3_119_728;
assign gate3_102_1478 = gate3_117_1453 & not_103_1477;
assign not_103_1477 = ~xor_109_1330;
assign gate3_98_1602 = gate3_88_1576 & not_99_1601;
assign not_99_1601 = ~gate3_85_1576;
assign gate3_85_1576 = not_86_1575 | not_121_1529;
assign not_121_1529 = ~xor_121_1528;
assign xor_121_1528 = gate3_104_728 ^ not_92_1504;
assign not_86_1575 = ~gate3_89_1555;
assign gate3_89_1555 = gate3_82_1503 | gate3_104_1528;
assign gate3_104_1528 = gate3_80_728 & not_85_1504;
assign gate3_82_1503 = not_114_1454 & not_83_1502;
assign not_83_1502 = ~gate3_92_1478;
assign gate3_88_1576 = gate3_92_1555 | xor_131_1528;
assign not_94_1655 = ~xor_94_1654;
assign xor_94_1654 = gate3_1_1628 ^ xor_15_1576;
assign gate3_22_1749 = gate3_23_1743 & gate3_77_1706;
assign gate3_77_1706 = gate3_131_1693 & gate3_97_1654;
assign gate3_97_1654 = gate3_110_1628 | gate3_79_1576;
assign gate3_110_1628 = gate3_110_1602 & not_111_1627;
assign not_111_1627 = ~gate3_102_1576;
assign gate3_102_1576 = not_121_1529 & not_103_1575;
assign not_103_1575 = ~gate3_89_1555;
assign gate3_110_1602 = gate3_85_1576 & not_111_1601;
assign not_111_1601 = ~xor_96_1576;
assign gate3_131_1693 = xor_4_1602 | gate3_1_1679;
assign gate3_23_1743 = gate3_23_1736 & not_24_1742;
assign not_24_1742 = ~gate3_97_1706;
assign gate3_97_1706 = gate3_1_1693 | gate3_137_1679;
assign gate3_137_1679 = gate3_108_1654 | gate3_111_1654;
assign gate3_111_1654 = gate3_132_1628 | not_112_1653;
assign not_112_1653 = ~gate3_135_1628;
assign gate3_135_1628 = gate3_132_1602 | gate3_102_1576;
assign gate3_132_1602 = gate3_88_1576 & not_133_1601;
assign not_133_1601 = ~gate3_99_1576;
assign gate3_132_1628 = xor_96_1576 & gate3_129_1602;
assign gate3_129_1602 = gate3_113_1576 | gate3_88_1576;
assign gate3_113_1576 = xor_145_1528 & not_114_1575;
assign not_114_1575 = ~gate3_99_1555;
assign xor_145_1528 = gate3_99_1503 ^ xor_143_1453;
assign xor_143_1453 = gate3_143_728 ^ not_147_1431;
assign not_147_1431 = ~xor_147_1430;
assign xor_147_1430 = not_148_1280 ^ gate3_133_1394;
assign gate3_133_1394 = gate3_133_1366 & gate3_129_1279;
assign gate3_129_1279 = xor_112_1182 | not_130_1278;
assign not_130_1278 = ~gate3_139_1233;
assign gate3_133_1366 = gate3_106_1330 | xor_135_1279;
assign not_148_1280 = ~xor_148_1279;
assign xor_148_1279 = gate3_147_1233 ^ gate3_90_983;
assign gate3_90_983 = gate3_124_857 & not_91_982;
assign not_91_982 = ~gate3_127_857;
assign gate3_127_857 = lever[38] & gate3_127_774;
assign gate3_127_774 = gate3_92_728 & gate3_128_728;
assign gate3_124_857 = gate3_140_728 | gate3_127_774;
assign gate3_140_728 = lever[19] & lever[38];
assign gate3_147_1233 = gate3_129_1108 | gate3_109_1182;
assign gate3_109_1182 = gate3_134_728 & not_110_1181;
assign not_110_1181 = ~not_139_1109;
assign gate3_129_1108 = gate3_145_1054 & gate3_151_774;
assign gate3_143_728 = lever[18] & lever[39];
assign gate3_99_1503 = gate3_126_1453 | gate3_106_1478;
assign gate3_106_1478 = gate3_131_728 & xor_133_1453;
assign gate3_126_1453 = gate3_133_1430 & xor_139_1366;
assign gate3_108_1654 = not_109_1653 & gate3_6_1628;
assign not_109_1653 = ~gate3_129_1628;
assign gate3_129_1628 = gate3_1_1602 & not_130_1627;
assign not_130_1627 = ~xor_17_1602;
assign gate3_23_1736 = gate3_21_1728 & not_24_1735;
assign not_24_1735 = ~not_122_1629;
assign not_122_1629 = ~xor_122_1628;
assign xor_122_1628 = xor_84_1602 ^ gate3_87_1602;
assign gate3_21_1728 = gate3_52_1654 & gate3_49_1720;
assign gate3_49_1720 = not_113_1603 & gate3_50_1714;
assign gate3_50_1714 = gate3_94_1706 & not_51_1713;
assign not_51_1713 = ~gate3_32_1602;
assign gate3_94_1706 = gate3_115_1628 & gate3_134_1693;
assign gate3_134_1693 = gate3_134_1679 & gate3_120_1602;
assign gate3_120_1602 = gate3_91_1576 | xor_145_1528;
assign gate3_91_1576 = not_111_1479 & not_92_1575;
assign not_92_1575 = ~gate3_99_1555;
assign gate3_134_1679 = not_135_1678 & gate3_105_1654;
assign gate3_105_1654 = gate3_108_1555 & gate3_118_1628;
assign gate3_118_1628 = gate3_123_1602 & not_119_1627;
assign not_119_1627 = ~gate3_115_1555;
assign gate3_115_1555 = gate3_129_1394 & gate3_142_1528;
assign gate3_142_1528 = xor_143_1453 | not_143_1527;
assign not_143_1527 = ~gate3_99_1503;
assign gate3_129_1394 = gate3_137_728 & gate3_150_1366;
assign gate3_150_1366 = gate3_121_1330 | gate3_116_1330;
assign gate3_116_1330 = gate3_139_1279 & not_117_1329;
assign not_117_1329 = ~gate3_129_1279;
assign gate3_139_1279 = gate3_147_1233 | gate3_90_983;
assign gate3_121_1330 = gate3_145_1279 | gate3_127_857;
assign gate3_145_1279 = gate3_147_1233 & gate3_90_983;
assign gate3_137_728 = lever[19] & lever[39];
assign gate3_123_1602 = gate3_123_1478 & gate3_110_1576;
assign gate3_110_1576 = not_111_1575 & gate3_118_1555;
assign gate3_118_1555 = gate3_148_1528 & not_119_1554;
assign not_119_1554 = ~gate3_40_1478;
assign gate3_148_1528 = gate3_154_1279 & gate3_113_1503;
assign gate3_113_1503 = gate3_145_1394 & gate3_131_1478;
assign gate3_131_1478 = gate3_150_1453 | gate3_177_1054;
assign gate3_177_1054 = gate3_115_983 | gate3_196_857;
assign gate3_196_857 = gate3_226_774 | gate3_260_728;
assign gate3_260_728 = lever[39] & not_261_727;
assign not_261_727 = ~lever[19];
assign gate3_226_774 = gate3_176_728 & not_227_773;
assign not_227_773 = ~xor_173_728;
assign xor_173_728 = lever[19] ^ lever[39];
assign gate3_176_728 = lever[38] & not_177_727;
assign not_177_727 = ~lever[18];
assign gate3_115_983 = gate3_193_857 & not_116_982;
assign not_116_982 = ~gate3_166_774;
assign gate3_166_774 = xor_173_728 | xor_179_728;
assign xor_179_728 = lever[18] ^ lever[38];
assign gate3_193_857 = gate3_257_728 | gate3_223_774;
assign gate3_223_774 = not_224_773 & gate3_185_728;
assign gate3_185_728 = lever[36] & not_186_727;
assign not_186_727 = ~lever[16];
assign not_224_773 = ~xor_182_728;
assign xor_182_728 = lever[17] ^ lever[37];
assign gate3_257_728 = lever[37] & not_258_727;
assign not_258_727 = ~lever[17];
assign gate3_150_1453 = gate3_93_983 & gate3_150_1430;
assign gate3_150_1430 = gate3_150_1394 | gate3_174_1054;
assign gate3_174_1054 = gate3_254_728 | gate3_112_983;
assign gate3_112_983 = gate3_190_857 & not_113_982;
assign not_113_982 = ~gate3_211_774;
assign gate3_211_774 = gate3_206_728 | xor_218_728;
assign xor_218_728 = lever[15] ^ lever[35];
assign gate3_206_728 = not_207_727 & lever[14];
assign not_207_727 = ~lever[34];
assign gate3_190_857 = gate3_205_774 | gate3_208_774;
assign gate3_208_774 = gate3_212_728 | gate3_251_728;
assign gate3_251_728 = lever[33] & not_252_727;
assign not_252_727 = ~lever[13];
assign gate3_212_728 = lever[34] & not_213_727;
assign not_213_727 = ~lever[14];
assign gate3_205_774 = gate3_209_728 & not_206_773;
assign not_206_773 = ~xor_215_728;
assign xor_215_728 = lever[33] ^ lever[13];
assign gate3_209_728 = lever[32] & not_210_727;
assign not_210_727 = ~lever[12];
assign gate3_254_728 = lever[35] & not_255_727;
assign not_255_727 = ~lever[15];
assign gate3_150_1394 = gate3_162_1054 & not_151_1393;
assign not_151_1393 = ~gate3_159_1366;
assign gate3_159_1366 = gate3_168_1054 & gate3_127_1330;
assign gate3_127_1330 = gate3_156_857 | gate3_158_1279;
assign gate3_158_1279 = gate3_158_1233 & gate3_180_857;
assign gate3_180_857 = gate3_242_728 & gate3_193_774;
assign gate3_193_774 = gate3_158_728 | xor_155_728;
assign xor_155_728 = lever[27] ^ lever[7];
assign gate3_158_728 = not_159_727 | lever[6];
assign not_159_727 = ~lever[26];
assign gate3_242_728 = not_243_727 | lever[7];
assign not_243_727 = ~lever[27];
assign gate3_158_1233 = gate3_160_774 | gate3_124_1182;
assign gate3_124_1182 = gate3_203_728 & gate3_145_1108;
assign gate3_145_1108 = gate3_165_1054 | gate3_172_774;
assign gate3_172_774 = gate3_197_728 | gate3_200_728;
assign gate3_200_728 = lever[4] & not_201_727;
assign not_201_727 = ~lever[24];
assign gate3_197_728 = not_198_727 & lever[5];
assign not_198_727 = ~lever[25];
assign gate3_165_1054 = gate3_99_983 & gate3_174_857;
assign gate3_174_857 = gate3_169_774 & gate3_190_774;
assign gate3_190_774 = gate3_164_728 | gate3_167_728;
assign gate3_167_728 = lever[2] | not_168_727;
assign not_168_727 = ~lever[22];
assign gate3_164_728 = not_165_727 & lever[3];
assign not_165_727 = ~lever[23];
assign gate3_169_774 = gate3_191_728 & gate3_194_728;
assign gate3_194_728 = lever[3] | not_195_727;
assign not_195_727 = ~lever[23];
assign gate3_191_728 = lever[4] | not_192_727;
assign not_192_727 = ~lever[24];
assign gate3_99_983 = gate3_168_857 | gate3_163_774;
assign gate3_163_774 = gate3_164_728 | xor_170_728;
assign xor_170_728 = lever[2] ^ lever[22];
assign gate3_168_857 = gate3_146_728 & gate3_157_774;
assign gate3_157_774 = xor_149_728 | gate3_152_728;
assign gate3_152_728 = lever[0] & not_153_727;
assign not_153_727 = ~lever[20];
assign xor_149_728 = lever[1] ^ lever[21];
assign gate3_146_728 = lever[1] | not_147_727;
assign not_147_727 = ~lever[21];
assign gate3_203_728 = lever[5] | not_204_727;
assign not_204_727 = ~lever[25];
assign gate3_160_774 = xor_161_728 | xor_155_728;
assign xor_161_728 = lever[26] ^ lever[6];
assign gate3_156_857 = gate3_178_774 | gate3_184_774;
assign gate3_184_774 = xor_236_728 | xor_239_728;
assign xor_239_728 = lever[29] ^ lever[9];
assign xor_236_728 = lever[8] ^ lever[28];
assign gate3_178_774 = xor_224_728 | xor_230_728;
assign xor_230_728 = lever[10] ^ lever[30];
assign xor_224_728 = lever[31] ^ lever[11];
assign gate3_168_1054 = gate3_109_983 & gate3_186_857;
assign gate3_186_857 = gate3_199_774 & gate3_248_728;
assign gate3_248_728 = lever[11] | not_249_727;
assign not_249_727 = ~lever[31];
assign gate3_199_774 = xor_224_728 | gate3_227_728;
assign gate3_227_728 = lever[10] | not_228_727;
assign not_228_727 = ~lever[30];
assign gate3_109_983 = gate3_178_774 | gate3_183_857;
assign gate3_183_857 = gate3_245_728 & gate3_196_774;
assign gate3_196_774 = gate3_233_728 | xor_239_728;
assign gate3_233_728 = lever[8] | not_234_727;
assign not_234_727 = ~lever[28];
assign gate3_245_728 = lever[9] | not_246_727;
assign not_246_727 = ~lever[29];
assign gate3_162_1054 = not_221_729 & not_163_1053;
assign not_163_1053 = ~gate3_96_983;
assign gate3_96_983 = xor_215_728 | gate3_145_857;
assign gate3_145_857 = xor_218_728 | gate3_175_774;
assign gate3_175_774 = gate3_206_728 | gate3_212_728;
assign not_221_729 = ~xor_221_728;
assign xor_221_728 = lever[12] ^ lever[32];
assign gate3_93_983 = not_188_729 & not_94_982;
assign not_94_982 = ~gate3_139_857;
assign gate3_139_857 = gate3_166_774 | xor_182_728;
assign not_188_729 = ~xor_188_728;
assign xor_188_728 = lever[16] ^ lever[36];
assign gate3_145_1394 = gate3_56_1366 | gate3_156_1366;
assign gate3_156_1366 = not_124_1331 & not_157_1365;
assign not_157_1365 = ~gate3_151_1279;
assign gate3_151_1279 = gate3_20_1182 | not_85_1234;
assign not_124_1331 = ~xor_124_1330;
assign xor_124_1330 = gate3_54_1233 ^ not_51_1280;
assign gate3_154_1279 = gate3_150_1233 & gate3_154_774;
assign gate3_154_774 = xor_149_728 & gate3_56_728;
assign gate3_150_1233 = gate3_98_1054 | gate3_121_1182;
assign gate3_121_1182 = not_57_1109 & not_85_858;
assign not_111_1575 = ~gate3_106_1503;
assign gate3_106_1503 = gate3_116_1478 & xor_141_1394;
assign xor_141_1394 = gate3_137_728 ^ gate3_150_1366;
assign gate3_116_1478 = gate3_138_1453 | not_117_1477;
assign not_117_1477 = ~gate3_136_1394;
assign gate3_136_1394 = gate3_133_1366 | not_148_1280;
assign gate3_138_1453 = gate3_143_728 & not_139_1452;
assign not_139_1452 = ~not_147_1431;
assign gate3_123_1478 = gate3_56_1366 | not_147_1454;
assign not_147_1454 = ~xor_147_1453;
assign xor_147_1453 = not_44_1430 ^ not_40_1431;
assign gate3_108_1555 = gate3_142_1528 | not_109_1554;
assign not_109_1554 = ~not_109_1504;
assign not_109_1504 = ~xor_109_1503;
assign xor_109_1503 = gate3_116_1478 ^ xor_141_1394;
assign not_135_1678 = ~gate3_125_1555;
assign gate3_125_1555 = gate3_26_1528 | not_126_1554;
assign not_126_1554 = ~gate3_29_1528;
assign gate3_115_1628 = not_116_1627 & gate3_136_1528;
assign gate3_136_1528 = gate3_23_1503 | xor_30_1503;
assign not_116_1627 = ~gate3_117_1602;
assign gate3_117_1602 = gate3_32_1528 | not_118_1601;
assign not_118_1601 = ~gate3_105_1576;
assign gate3_105_1576 = gate3_129_1394 | gate3_102_1555;
assign gate3_102_1555 = gate3_142_1528 & not_109_1504;
assign not_113_1603 = ~xor_113_1602;
assign xor_113_1602 = not_10_1556 ^ gate3_18_1576;
assign gate3_20_1743 = gate3_79_1654 | gate3_20_1736;
assign gate3_20_1736 = gate3_28_1628 & not_21_1735;
assign not_21_1735 = ~gate3_1_1728;
assign gate3_79_1654 = gate3_34_1628 & not_80_1653;
assign not_80_1653 = ~xor_41_1628;
assign gate3_18_1764 = xor_41_1628 | not_19_1763;
assign not_19_1763 = ~gate3_1_1756;
assign not_10_1799 = ~gate3_9_1793;
assign gate3_9_1793 = xor_11_1679 & gate3_1_1785;
assign not_4_1814 = ~xor_4_1813;
assign xor_4_1813 = xor_54_1679 ^ gate3_1_1805;
assign not_9_1828 = ~xor_9_1827;
assign xor_9_1827 = xor_64_1679 ^ gate3_1_1819;
assign gate3_9_1849 = xor_86_1679 | gate3_6_1841;
assign not_5_1891 = ~gate3_4_1876;
assign gate3_4_1876 = gate3_75_1654 & not_5_1875;
assign not_5_1875 = ~gate3_6_1866;
assign gate3_7_1901 = gate3_1_1892 | xor_90_1602;
assign gate3_1_1929 = gate3_1_1922 | xor_82_1576;
assign gate3_1_1922 = gate3_1_1915 & gate3_73_1576;

cover property(lamp_1_1938);

endmodule
